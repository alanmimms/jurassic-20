module cha27(
      input  cam_sel_1_h                       /* <br1> */,
      input  cam_sel_2_h                       /* <bs1> */,
      input  con_wr_even_par_dir_l             /* <ad2> */,
      output csh_0_any_wr_l                    /* <al2> */,
      input  csh_0_wr_en_l                     /* <al1> */,
      output csh_1_any_wr_l                    /* <aj2> */,
      input  csh_1_wr_en_l                     /* <am1> */,
      output csh_2_any_wr_l                    /* <bl2> */,
      input  csh_2_wr_en_l                     /* <aj1> */,
      output csh_3_any_wr_l                    /* <be2> */,
      input  csh_3_wr_en_l                     /* <ak2> */,
      input  csh_adr_wr_pulse_l                /* <bj2> */,
      output csh_dir_14_0_h                    /* <da1> */,
      output csh_dir_14_1_h                    /* <cj1> */,
      output csh_dir_14_2_h                    /* <dl2> */,
      output csh_dir_14_3_h                    /* <df2> */,
      output csh_dir_15_0_h                    /* <cm1> */,
      output csh_dir_15_1_h                    /* <cd1> */,
      output csh_dir_15_2_h                    /* <dl1> */,
      output csh_dir_15_3_h                    /* <de1> */,
      output csh_dir_16_0_h                    /* <cl1> */,
      output csh_dir_16_1_h                    /* <cc1> */,
      output csh_dir_16_2_h                    /* <ca1> */,
      output csh_dir_16_3_h                    /* <dc1> */,
      output csh_dir_17_0_h                    /* <cp1> */,
      output csh_dir_17_1_h                    /* <cf1> */,
      output csh_dir_17_2_h                    /* <ce1> */,
      output csh_dir_17_3_h                    /* <dd2> */,
      output csh_dir_18_0_h                    /* <dr1> */,
      output csh_dir_18_1_h                    /* <dt2> */,
      output csh_dir_18_2_h                    /* <ef1> */,
      output csh_dir_18_3_h                    /* <ea1> */,
      output csh_dir_19_0_h                    /* <dn1> */,
      output csh_dir_19_1_h                    /* <ds1> */,
      output csh_dir_19_2_h                    /* <ee2> */,
      output csh_dir_19_3_h                    /* <ec1> */,
      output csh_dir_20_0_h                    /* <dj1> */,
      output csh_dir_20_1_h                    /* <dm1> */,
      output csh_dir_20_2_h                    /* <du2> */,
      output csh_dir_20_3_h                    /* <dr2> */,
      output csh_dir_21_0_h                    /* <dk1> */,
      output csh_dir_21_1_h                    /* <dm2> */,
      output csh_dir_21_2_h                    /* <dv2> */,
      output csh_dir_21_3_h                    /* <ds2> */,
      output csh_dir_22_0_h                    /* <eh2> */,
      output csh_dir_22_1_h                    /* <ep2> */,
      output csh_dir_22_2_h                    /* <fd1> */,
      output csh_dir_22_3_h                    /* <es2> */,
      output csh_dir_23_0_h                    /* <ef2> */,
      output csh_dir_23_1_h                    /* <ep1> */,
      output csh_dir_23_2_h                    /* <fe1> */,
      output csh_dir_23_3_h                    /* <er1> */,
      output csh_dir_24_0_h                    /* <ed1> */,
      output csh_dir_24_1_h                    /* <ek2> */,
      output csh_dir_24_2_h                    /* <eu2> */,
      output csh_dir_24_3_h                    /* <el2> */,
      output csh_dir_25_0_h                    /* <ee1> */,
      output csh_dir_25_1_h                    /* <el1> */,
      output csh_dir_25_2_h                    /* <ev2> */,
      output csh_dir_25_3_h                    /* <em1> */,
      output csh_dir_26_0_h                    /* <fd2> */,
      output csh_dir_26_1_h                    /* <fl2> */,
      output csh_dir_26_2_h                    /* <fu2> */,
      output csh_dir_26_3_h                    /* <fk1> */,
      output csh_dir_par_0_h                   /* <fr2> */,
      output csh_dir_par_1_h                   /* <fp1> */,
      output csh_dir_par_2_h                   /* <fn1> */,
      output csh_dir_par_3_h                   /* <fp2> */,
      output csh_wd_0_wr_h                     /* <au2> */,
      output csh_wd_1_wr_h                     /* <am2> */,
      output csh_wd_2_wr_h                     /* <bd2> */,
      output csh_wd_3_wr_h                     /* <av2> */,
      input  csh_wr_out_en_l                   /* <ar2> */,
      input  csh_wr_sel_all_h                  /* <as2> */,
      input  csh_wr_wd_0_en_h                  /* <ae1> */,
      input  csh_wr_wd_1_en_h                  /* <af1> */,
      input  csh_wr_wd_2_en_h                  /* <aa1> */,
      input  csh_wr_wd_3_en_h                  /* <ad1> */,
      input  csh_wr_wr_data_h                  /* <af2> */,
      input  csh_wr_wr_pulse_l                 /* <bf2> */,
      input  mbx_csh_adr_27_h                  /* <as1> */,
      input  mbx_csh_adr_28_h                  /* <an1> */,
      input  mbx_csh_adr_29_h                  /* <be1> */,
      input  mbx_csh_adr_30_h                  /* <ba1> */,
      input  mbx_csh_adr_31_h                  /* <bp1> */,
      input  mbx_csh_adr_32_h                  /* <bl1> */,
      input  mbx_csh_adr_33_h                  /* <bf1> */,
      input  pma_14_h                          /* <cv2> */,
      input  pma_14to26_par_h                  /* <ae2> */,
      input  pma_15_h                          /* <cu2> */,
      input  pma_16_h                          /* <cd2> */,
      input  pma_17_h                          /* <cl2> */,
      input  pma_18_h                          /* <df1> */,
      input  pma_19_h                          /* <dp1> */,
      input  pma_20_h                          /* <ed2> */,
      input  pma_21_h                          /* <ej1> */,
      input  pma_22_h                          /* <fj1> */,
      input  pma_23_h                          /* <fa1> */,
      input  pma_24_h                          /* <ek1> */,
      input  pma_25_h                          /* <es1> */,
      input  pma_26_h                          /* <dd1> */,
      input  vma_27_g_h                        /* <ar1> */,
      input  vma_28_g_h                        /* <ap1> */,
      input  vma_29_g_h                        /* <bd1> */,
      input  vma_30_g_h                        /* <bc1> */,
      input  vma_31_g_h                        /* <bm2> */,
      input  vma_32_g_h                        /* <bm1> */,
      input  vma_33_g_h                        /* <bj1> */
);

`include "cha27nets.svh"

endmodule	// cha27
