module ctl36(
      input  apr2_clk_c_h                      /* <aa1> */,
      input  apr3_coni_or_datai_l              /* <el1> */,
      input  apr3_cono_or_datao_h              /* <ba1> */,
      input  apr_ebus_return_h                 /* <an1> */,
      input  ar_00_c_h                         /* <er1> */,
      input  arx_18_b_h                        /* <fk2> */,
      input  clk4_resp_mbox_h                  /* <fl2> */,
      input  clk_resp_sim_h                    /* <fk1> */,
      input  clk_sbr_call_h                    /* <af1> */,
      input  con_condSldiag_func_l             /* <dd1> */,
      input  con_cond_en_00to07_l              /* <bc1> */,
      input  con_fm_xfer_h                     /* <fv2> */,
      input  con_pcPl1_inh_h                   /* <es2> */,
      input  con_pi_cycle_b_h                  /* <bh2> */,
      input  cra3_disp_00_h                    /* <et2> */,
      input  cra3_disp_01_h                    /* <es1> */,
      input  cra3_disp_02_h                    /* <df2> */,
      input  cra3_disp_03_h                    /* <de2> */,
      input  cra3_disp_04_h                    /* <dj2> */,
      input  cram_Nr_00_c_h                    /* <er2> */,
      input  cram_Nr_01_c_h                    /* <ep1> */,
      input  cram_Nr_02_c_h                    /* <dp1> */,
      input  cram_Nr_03_c_h                    /* <dr1> */,
      input  cram_Nr_04_c_h                    /* <ek2> */,
      input  cram_Nr_05_c_h                    /* <dp2> */,
      input  cram_Nr_06_c_h                    /* <en1> */,
      input  cram_Nr_07_c_h                    /* <dl1> */,
      input  cram_Nr_08_c_h                    /* <bm1> */,
      input  cram_ad_cry_h                     /* <bd2> */,
      input  cram_arm_sel_1_h                  /* <fh2> */,
      input  cram_arm_sel_2_h                  /* <ev2> */,
      input  cram_arm_sel_4_h                  /* <em1> */,
      input  cram_arxm_sel_1_h                 /* <ft2> */,
      input  cram_arxm_sel_2_h                 /* <fm2> */,
      input  cram_arxm_sel_4_h                 /* <eu2> */,
      input  cram_cond_03_a_l                  /* <bd1> */,
      input  cram_cond_04_a_l                  /* <be1> */,
      input  cram_cond_05_a_l                  /* <bf2> */,
      input  cram_mq_sel_h                     /* <ff1> */,
      output ctl1_condSlarGETSexp_h            /* <dc1> */,
      output ctl1_disp_ret_l                   /* <cs2> */,
      output ctl1_load_pc_l                    /* <cp2> */,
      output ctl1_specSlclr_fpd_h              /* <cm1> */,
      output ctl1_specSlflag_ctl_h             /* <ck2> */,
      output ctl1_specSlscm_alt_h              /* <cl2> */,
      output ctl1_specSlsp_mem_cycle_h         /* <cl1> */,
      output ctl1_spec_mtr_ctl_l               /* <da1> */,
      output ctl2_ebus_xfer_h                  /* <dd2> */,
      output ctl2_spec_call_l                  /* <em2> */,
      output ctl3_diag_clk_edp_h               /* <be2> */,
      output ctl3_diag_ctl_func_00x_l          /* <at2> */,
      output ctl3_diag_diag_04_h               /* <fm1> */,
      output ctl3_diag_diag_04_l               /* <fn1> */,
      output ctl3_diag_force_extend_h          /* <fr1> */,
      output ctl3_diag_force_extend_l          /* <fr2> */,
      output ctl3_diag_ld_ebus_reg_h           /* <fp1> */,
      output ctl3_diag_ld_ebus_reg_l           /* <df1> */,
      output ctl3_diag_ld_func_04x_l           /* <ap2> */,
      output ctl3_diag_ld_func_072_l           /* <aj1> */,
      output ctl3_diag_ld_func_073_l           /* <af2> */,
      output ctl3_diag_ld_func_075_l           /* <ad2> */,
      output ctl3_diag_rd_func_11x_l           /* <ck1> */,
      output ctl3_diag_spare_h                 /* <fj1> */,
      input  ctl3_diag_spare_l                 /* <fj2> */,
      output ctl3_diag_sync_func_074_l         /* <ae1> */,
      output ctl_ad_long_h                     /* <bl2> */,
      output ctl_ad_to_ebus_l_h                /* <br1> */,
      output ctl_ad_to_ebus_r_h                /* <br2> */,
      output ctl_adx_cry_36_a_h                /* <bs2> */,
      output ctl_adx_cry_36_h                  /* <bt2> */,
      output ctl_ar_00to08_load_l              /* <dm1> */,
      output ctl_ar_00to11_clr_h               /* <ef1> */,
      output ctl_ar_09to17_load_l              /* <ee2> */,
      output ctl_ar_12to17_clr_h               /* <ej1> */,
      output ctl_arl_sel_1_h                   /* <ee1> */,
      output ctl_arl_sel_2_h                   /* <ec1> */,
      output ctl_arl_sel_4_h                   /* <ed2> */,
      output ctl_arr_clr_h                     /* <ej2> */,
      output ctl_arr_load_a_l                  /* <ed1> */,
      output ctl_arr_load_b_l                  /* <dk2> */,
      output ctl_arr_sel_1_h                   /* <ef2> */,
      output ctl_arr_sel_2_h                   /* <ea1> */,
      output ctl_arx_load_h                    /* <dn1> */,
      output ctl_arxl_sel_1_h                  /* <fc1> */,
      output ctl_arxl_sel_2_h                  /* <fd2> */,
      output ctl_arxr_sel_1_h                  /* <fa1> */,
      output ctl_arxr_sel_2_h                  /* <fd1> */,
      output ctl_console_control_h             /* <dj1> */,
      output ctl_dispSlnicond_h                /* <bj1> */,
      output ctl_ebus_e_to_t_en_h              /* <am1> */,
      output ctl_ebus_parity_out_e_h           /* <bm2> */,
      output ctl_ebus_t_to_e_en_h              /* <bk1> */,
      output ctl_ebus_xfer_l                   /* <de1> */,
      output ctl_gen_cry_18_h                  /* <cm2> */,
      output ctl_inh_cry_18_l                  /* <bl1> */,
      output ctl_mq_sel_1_h                    /* <bu2> */,
      output ctl_mq_sel_2_h                    /* <bv2> */,
      output ctl_mqm_en_h                      /* <dh2> */,
      output ctl_mqm_sel_1_h                   /* <dl2> */,
      output ctl_mqm_sel_2_h                   /* <dk1> */,
      output ctl_specSlflag_ctl_l              /* <cu2> */,
      output ctl_specSlgen_cry_18_h            /* <aa2> */,
      output ctl_specSlsave_flags_l            /* <cr2> */,
      output diag_04_a_h                       /* <bp2> */,
      output diag_04_a_l                       /* <fe1> */,
      output diag_04_b_h                       /* <as2> */,
      output diag_04_b_l                       /* <as1> */,
      output diag_05_a_h                       /* <bp1> */,
      output diag_05_a_l                       /* <fe2> */,
      output diag_05_b_h                       /* <al2> */,
      output diag_05_b_l                       /* <al1> */,
      output diag_06_a_h                       /* <cr1> */,
      output diag_06_a_l                       /* <ff2> */,
      output diag_06_b_h                       /* <am2> */,
      output diag_06_b_l                       /* <ak2> */,
      output diag_channel_clk_stop_h           /* <fp2> */,
      output diag_control_func_01x_l           /* <av2> */,
      output diag_load_func_05x_l              /* <ap1> */,
      output diag_load_func_06x_l              /* <ar1> */,
      output diag_load_func_070_l              /* <ak1> */,
      output diag_load_func_071_l              /* <ah2> */,
      output diag_mem_reset_h                  /* <bs1> */,
      output diag_read_func_10x_l              /* <cj2> */,
      output diag_read_func_12x_h              /* <bf1> */,
      output diag_read_func_13x_l              /* <ch2> */,
      output diag_read_func_14x_l              /* <cj1> */,
      output diag_read_func_15x_l              /* <cf2> */,
      output diag_read_func_16x_l              /* <ce1> */,
      output diag_read_func_17x_l              /* <cf1> */,
      output ebus_d24_e_h                      /* <dr2> */,
      output ebus_d25_e_h                      /* <ds1> */,
      output ebus_d26_e_h                      /* <ds2> */,
      output ebus_d27_e_h                      /* <dt2> */,
      output ebus_d28_e_h                      /* <du2> */,
      input  ebus_ds00_e_h                     /* <ce2> */,
      input  ebus_ds01_e_h                     /* <cd2> */,
      input  ebus_ds02_e_h                     /* <cd1> */,
      input  ebus_ds03_e_h                     /* <cc1> */,
      input  ebus_ds04_e_h                     /* <ca1> */,
      input  ebus_ds05_e_h                     /* <ae2> */,
      input  ebus_ds06_e_h                     /* <aj2> */,
      input  ebus_ds_strobe_e_h                /* <bj2> */,
      input  mcl1_memSlarl_ind_h               /* <ac1> */,
      input  mcl4_short_stack_h                /* <cn1> */,
      input  mcl5_18_bit_ea_h                  /* <fs2> */,
      input  mcl5_23_bit_ea_h                  /* <fs1> */,
      input  mcl_load_ar_h                     /* <fl1> */,
      input  mcl_load_arx_h                    /* <fu2> */,
      input  mr_reset_04_h                     /* <ep2> */,
      input  pi5_gate_ttl_to_ecl_l             /* <el2> */,
      input  shm1_ar_par_odd_a_l               /* <bk2> */
);

`include "ctl36nets.svh"

endmodule	// ctl36
