module delay_line(input bit in, output bit out);
  always_comb out = in;
endmodule // delay_line
