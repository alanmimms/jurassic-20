module top(input clk);

   

endmodule // top
