module edp43(
      input  ad_16_h                           /* <cp2> */,
      input  ad_17_h                           /* <el2> */,
      output ad_18_a_h                         /* <ck1> */,
      output ad_18_a_l                         /* <cn1> */,
      output ad_18_h                           /* <ep2> */,
      output ad_18to23Eq0_l                    /* <at2> */,
      output ad_19_h                           /* <dl1> */,
      output ad_20_h                           /* <dr2> */,
      output ad_21_h                           /* <dr1> */,
      output ad_22_a_h                         /* <cf2> */,
      output ad_22_h                           /* <cp1> */,
      output ad_23_a_h                         /* <ce1> */,
      output ad_23_h                           /* <el1> */,
      input  ad_24_h                           /* <ep1> */,
      output ad_cg_18_h                        /* <am1> */,
      output ad_cg_20_h                        /* <am2> */,
      output ad_cp_18_h                        /* <aj1> */,
      output ad_cp_20_h                        /* <af1> */,
      output ad_cry_19_h                       /* <cu2> */,
      output ad_cry_19_l                       /* <ct2> */,
      input  ad_cry_24_h                       /* <al1> */,
      output ad_ex_16_h                        /* <cv2> */,
      output ad_ex_17_h                        /* <cr1> */,
      output ad_overflow_18_l                  /* <cl2> */,
      input  adx_17_h                          /* <es2> */,
      output adx_18_a_h                        /* <cf1> */,
      output adx_18_h                          /* <cj2> */,
      output adx_22_h                          /* <dk1> */,
      output adx_23_h                          /* <es1> */,
      input  adx_24_h                          /* <cj1> */,
      output adx_cg_18_h                       /* <al2> */,
      output adx_cg_21_h                       /* <ak2> */,
      output adx_cp_18_h                       /* <ae1> */,
      output adx_cp_21_h                       /* <af2> */,
      input  adx_cry_24_h                      /* <ak1> */,
      input  apr_fm_adr_10_h                   /* <fr2> */,
      input  apr_fm_adr_1_h                    /* <fp2> */,
      input  apr_fm_adr_2_h                    /* <fs1> */,
      input  apr_fm_adr_4_h                    /* <fn1> */,
      input  apr_fm_block_1_h                  /* <fr1> */,
      input  apr_fm_block_2_h                  /* <fm1> */,
      input  apr_fm_block_4_h                  /* <fp1> */,
      output ar_18_a_h                         /* <fj2> */,
      output ar_18_b_h                         /* <ft2> */,
      output ar_18_c_h                         /* <fs2> */,
      output ar_18_d_h                         /* <dm2> */,
      output ar_18_h                           /* <bk2> */,
      output ar_19_a_h                         /* <fc1> */,
      output ar_19_b_h                         /* <fu2> */,
      output ar_19_c_h                         /* <fv2> */,
      output ar_19_h                           /* <bl2> */,
      output ar_20_a_h                         /* <ff2> */,
      output ar_20_b_h                         /* <cl1> */,
      output ar_20_c_h                         /* <ch2> */,
      output ar_21_a_h                         /* <eu2> */,
      output ar_21_b_h                         /* <ck2> */,
      output ar_21_c_h                         /* <cm1> */,
      output ar_22_a_h                         /* <ev2> */,
      output ar_22_b_h                         /* <fk1> */,
      output ar_22_c_h                         /* <fk2> */,
      output ar_23_a_h                         /* <et2> */,
      output ar_23_b_h                         /* <fl2> */,
      output ar_23_c_h                         /* <fl1> */,
      input  ar_24_h                           /* <bk1> */,
      input  ar_25_h                           /* <bl1> */,
      input  armm_18_h                         /* <em2> */,
      input  armm_19_h                         /* <ea1> */,
      input  armm_20_h                         /* <ee1> */,
      input  armm_21_h                         /* <dd2> */,
      input  armm_22_h                         /* <de1> */,
      input  armm_23_h                         /* <ef2> */,
      output arx_18_a_h                        /* <as2> */,
      output arx_18_b_h                        /* <br2> */,
      output arx_18_h                          /* <ej2> */,
      output arx_19_a_h                        /* <as1> */,
      output arx_19_b_h                        /* <cm2> */,
      output arx_19_h                          /* <bd2> */,
      output arx_20_h                          /* <dc1> */,
      output arx_21_h                          /* <aj2> */,
      output arx_22_h                          /* <ac1> */,
      output arx_23_h                          /* <aa1> */,
      input  arx_24_h                          /* <ej1> */,
      input  arx_25_h                          /* <bd1> */,
      output br_18_a_h                         /* <bm2> */,
      input  br_24_a_h                         /* <bm1> */,
      output brx_18_h                          /* <be2> */,
      input  brx_24_h                          /* <be1> */,
      input  cache_data_18_b_h                 /* <em1> */,
      input  cache_data_19_b_h                 /* <ed2> */,
      input  cache_data_20_b_h                 /* <ee2> */,
      input  cache_data_21_b_h                 /* <dd1> */,
      input  cache_data_22_b_h                 /* <dl2> */,
      input  cache_data_23_b_h                 /* <cc1> */,
      input  clk_edp_18_h                      /* <cr2> */,
      input  con_fm_write_18to35_l             /* <ce2> */,
      input  cram_Nr_18_h                      /* <ar1> */,
      input  cram_Nr_19_h                      /* <ap1> */,
      input  cram_Nr_20_h                      /* <ba1> */,
      input  cram_Nr_21_h                      /* <ap2> */,
      input  cram_Nr_22_h                      /* <av2> */,
      input  cram_Nr_23_h                      /* <au2> */,
      input  cram_ad_boole_18_h                /* <an1> */,
      input  cram_ad_sel_1_18_h                /* <ad2> */,
      input  cram_ad_sel_2_18_h                /* <ah2> */,
      input  cram_ad_sel_4_18_h                /* <ae2> */,
      input  cram_ad_sel_8_18_h                /* <ad1> */,
      input  cram_ada_dis_18_h                 /* <bn1> */,
      input  cram_ada_sel_1_18_h               /* <bj1> */,
      input  cram_ada_sel_2_18_h               /* <bf2> */,
      input  cram_adb_sel_1_18_h               /* <bt2> */,
      input  cram_adb_sel_2_18_h               /* <bs1> */,
      input  cram_arm_sel_4_a_h                /* <er1> */,
      input  cram_arxm_sel_4_06_h              /* <ff1> */,
      input  cram_br_load_a_h                  /* <dj2> */,
      input  cram_brx_load_a_h                 /* <ar2> */,
      input  ctl_ad_to_ebus_r_h                /* <fe2> */,
      input  ctl_arr_clr_h                     /* <eh2> */,
      input  ctl_arr_load_a_l                  /* <ek2> */,
      input  ctl_arr_load_b_l                  /* <dh2> */,
      input  ctl_arr_sel_1_h                   /* <en1> */,
      input  ctl_arr_sel_2_h                   /* <ek1> */,
      input  ctl_arx_load_h                    /* <br1> */,
      input  ctl_arxr_sel_1_h                  /* <fj1> */,
      input  ctl_arxr_sel_2_h                  /* <fd2> */,
      input  ctl_mq_sel_1_h                    /* <bu2> */,
      input  ctl_mq_sel_2_h                    /* <bv2> */,
      input  ctl_mqm_en_h                      /* <dn1> */,
      input  ctl_mqm_sel_1_h                   /* <dj1> */,
      input  ctl_mqm_sel_2_h                   /* <dm1> */,
      input  diag_04_a_h                       /* <fd1> */,
      input  diag_05_a_h                       /* <fa1> */,
      input  diag_06_a_h                       /* <fe1> */,
      input  diag_read_func_12x_h              /* <ef1> */,
      output ebus_d18_e_h                      /* <dv2> */,
      output ebus_d19_e_h                      /* <ds2> */,
      output ebus_d20_e_h                      /* <dt2> */,
      output ebus_d21_e_h                      /* <dp1> */,
      output ebus_d22_e_h                      /* <dp2> */,
      output ebus_d23_e_h                      /* <du2> */,
      output edp_fm_parity_18to23_h            /* <fm2> */,
      input  mq_16_h                           /* <cs2> */,
      output mq_18_h                           /* <cd2> */,
      output mq_22_h                           /* <cs1> */,
      output mq_23_h                           /* <df1> */,
      input  mq_24_h                           /* <cd1> */,
      input  sh_18_h                           /* <ed1> */,
      input  sh_19_h                           /* <ec1> */,
      input  sh_20_h                           /* <ds1> */,
      input  sh_21_h                           /* <da1> */,
      input  sh_22_h                           /* <de2> */,
      input  sh_23_h                           /* <ca1> */,
      input  vma_held_or_pc_18_h               /* <bj2> */,
      input  vma_held_or_pc_19_h               /* <bh2> */,
      input  vma_held_or_pc_20_h               /* <bf1> */,
      input  vma_held_or_pc_21_h               /* <bp2> */,
      input  vma_held_or_pc_22_h               /* <bp1> */,
      input  vma_held_or_pc_23_h               /* <bc1> */
);

`include "edp43nets.svh"

endmodule	// edp43
