module wire6(input bit a, output bit q1, q2, q3, q4, q5, q6);
  always_comb begin
    q1 = a;
    q2 = a;
    q3 = a;
    q4 = a;
    q5 = a;
    q6 = a;
  end
endmodule // wire6
