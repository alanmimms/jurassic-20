module ctl;
`include "ctl.svh"
endmodule	// ctl
