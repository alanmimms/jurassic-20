module csh;
`include "csh.svh"
endmodule	// csh
