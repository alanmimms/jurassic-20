module chc;
`include "chc.svh"
endmodule	// chc
