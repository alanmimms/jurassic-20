module crm;
`include "crm.svh"
endmodule	// crm
