module mbx21(
  /* <er1> */  input ackn_pulse_l,
  /* <em1> */  input apr2_c_dir_p_err_h,
  /* <fd1> */  input apr6_ebox_cca_h,
  /* <dn1> */  input apr_ebox_sbus_diag_l,
  /* <dj2> */  input cache_exists_l,
  /* <ck2> */ output cache_to_mb_t4_l,
  /* <ej1> */  input ccl_ch_load_mb_l,
  /* <ah2> */  input ccl_ch_mb_sel_1_h,
  /* <ak2> */  input ccl_ch_mb_sel_2_h,
  /* <ds1> */  input ccl_chan_to_mem_h,
  /* <cp1> */  input ccw_cha_34_h,
  /* <br1> */  input ccw_cha_35_h,
  /* <an1> */  input ccw_wd0_req_h,
  /* <ap2> */  input ccw_wd1_req_h,
  /* <cn1> */  input ccw_wd2_req_h,
  /* <cl2> */  input ccw_wd3_req_h,
  /* <ej2> */  input chan_read_l,
  /* <cr2> */  input clk1_mbx_h,
  /* <es1> */  input con_cache_look_en_l,
  /* <ea1> */  input core_busy_a_h,
  /* <ef1> */  input core_rd_in_prog_h,
  /* <eh2> */  input csh1_cca_cyc_l,
  /* <dl1> */  input csh1_mb_cyc_l,
  /* <fs1> */  input csh1_mb_req_grant_l,
  /* <dk1> */  input csh1_pgrf_cyc_a_l,
  /* <fc1> */  input csh1_ready_to_go_h,
  /* <fs2> */  input csh1_ready_to_go_l,
  /* <dm2> */  input csh2_e_cache_wr_cyc_h,
  /* <cj2> */  input csh2_e_core_rd_rq_l,
  /* <cp2> */  input csh2_one_word_rd_l,
  /* <dr1> */  input csh3_adr_ready_l,
  /* <fp2> */  input csh3_any_val_hold_in_h,
  /* <fp1> */  input csh3_mb_wr_rq_clr_nxt_l,
  /* <el1> */  input csh4_one_word_wr_t0_l,
  /* <dl2> */  input csh4_writeback_t1_a_l,
  /* <ec1> */  input csh5_chan_t4_l,
  /* <ed2> */  input csh5_page_refill_t8_l,
  /* <ed1> */  input csh5_t2_l,
  /* <ev2> */  input csh6_cca_cyc_done_l,
  /* <eu2> */  input csh6_cca_inval_t4_l,
  /* <ep1> */  input csh6_ebox_load_reg_h,
  /* <dp1> */  input csh_adr_par_bad_l,
  /* <el2> */ output csh_chan_cyc_a_h,
  /* <du2> */  input csh_chan_cyc_l,
  /* <fd2> */  input csh_wd_0_val_h,
  /* <ad2> */  input csh_wd_0_wr_h,
  /* <er2> */  input csh_wd_1_val_h,
  /* <ac1> */  input csh_wd_1_wr_h,
  /* <fe2> */  input csh_wd_2_val_h,
  /* <ad1> */  input csh_wd_2_wr_h,
  /* <fj2> */  input csh_wd_3_val_h,
  /* <aa1> */  input csh_wd_3_wr_h,
  /* <dv2> */ output csh_wr_out_en_l,
  /* <cu2> */ output csh_wr_wd_0_en_h,
  /* <cs1> */ output csh_wr_wd_1_en_h,
  /* <ba1> */ output csh_wr_wd_2_en_h,
  /* <av2> */ output csh_wr_wd_3_en_h,
  /* <bn1> */  input diag_04_b_h,
  /* <bp1> */  input diag_05_b_h,
  /* <bl1> */  input diag_06_b_h,
  /* <dh2> */  input diag_load_func_071_l,
  /* <bk2> */  input diag_read_func_17x_l,
  /* <da1> */ output ebus_d30_e_h,
  /* <dc1> */ output ebus_d31_e_h,
  /* <dd2> */ output ebus_d32_e_h,
  /* <df2> */ output ebus_d33_e_h,
  /* <cc1> */ output ebus_d34_e_h,
  /* <ca1> */ output ebus_d35_e_h,
  /* <au2> */ output force_no_match_h,
  /* <fh2> */  input ir_ac_10_h,
  /* <ff2> */  input ir_ac_11_h,
  /* <ff1> */  input ir_ac_12_h,
  /* <bl2> */ output mb0_hold_in_h,
  /* <bm1> */ output mb1_hold_in_h,
  /* <bk1> */ output mb2_hold_in_h,
  /* <bj2> */ output mb3_hold_in_h,
  /* <as2> */ output mb_data_code_1_h,
  /* <as1> */ output mb_data_code_2_h,
  /* <ek2> */  input mb_in_sel_1_h,
  /* <ch2> */  input mb_in_sel_2_h,
  /* <cf1> */  input mb_in_sel_4_h,
  /* <am2> */  input mb_par_bit_in_h,
  /* <ar2> */ output mb_par_h,
  /* <ar1> */ output mb_req_hold_h,
  /* <ak1> */ output mb_sel_1_en_h,
  /* <cf2> */ output mb_sel_1_h,
  /* <ae1> */ output mb_sel_2_en_h,
  /* <bp2> */ output mb_sel_2_h,
  /* <af1> */ output mb_sel_hold_h,
  /* <ft2> */  input mbc2_csh_data_clr_t3_l,
  /* <ds2> */  input mbc3_a_change_coming_a_l,
  /* <al1> */  input mbc3_csh_wr_wr_data_l,
  /* <es2> */  input mbc3_inh_1st_mb_req_h,
  /* <bh2> */  input mbc4_core_adr_34_h,
  /* <bj1> */  input mbc4_core_adr_35_h,
  /* <ep2> */  input mbc4_core_data_val_Ng2_l,
  /* <ef2> */  input mbc4_mem_start_l,
  /* <de2> */ output mbx1_cache_bit_h,
  /* <fj1> */ output mbx1_cache_bit_l,
  /* <cm2> */ output mbx1_cca_all_pages_cyc_h,
  /* <fv2> */ output mbx1_cca_all_pages_cyc_l,
  /* <et2> */ output mbx1_cca_inval_t4_a_h,
  /* <df1> */ output mbx1_cca_req_l,
  /* <de1> */ output mbx1_cca_sel_1_h,
  /* <dd1> */ output mbx1_cca_sel_2_h,
  /* <cv2> */ output mbx1_csh_cca_inval_csh_h,
  /* <ct2> */ output mbx1_csh_cca_val_core_h,
  /* <fm1> */ output mbx1_csh_cca_val_core_l,
  /* <ap1> */ output mbx1_ebox_load_reg_h,
  /* <fu2> */ output mbx1_force_match_en_l,
  /* <fn1> */ output mbx1_refill_adr_en_h,
  /* <fr2> */ output mbx1_refill_adr_en_nxt_h,
  /* <fl2> */ output mbx2_cache_to_mb_34_h,
  /* <fe1> */ output mbx2_cache_to_mb_35_h,
  /* <dj1> */ output mbx2_chan_wr_cyc_l,
  /* <am1> */ output mbx2_mb_sel_hold_ff_h,
  /* <ee2> */ output mbx2_mb_sel_hold_l,
  /* <bs2> */ output mbx3_refill_hold_h,
  /* <bd1> */ output mbx3_sbus_diag_3_l,
  /* <ek1> */ output mbx4_cache_to_mb_done_l,
  /* <dk2> */ output mbx4_cache_to_mb_t2_l,
  /* <cm1> */ output mbx4_cache_to_mb_t4_a_l,
  /* <dt2> */ output mbx4_writeback_t2_h,
  /* <bc1> */ output mbx4_writeback_t2_l,
  /* <en1> */ output mbx5_csh_adr_par_err_l,
  /* <ce1> */ output mbx5_mb_req_in_h,
  /* <cd2> */ output mbx5_mem_rd_rq_in_h,
  /* <cd1> */ output mbx5_mem_to_c_en_l,
  /* <bt2> */ output mbx5_mem_wr_rq_in_h,
  /* <cs2> */ output mbx5_mem_wr_rq_in_l,
  /* <bs1> */ output mbx5_rq_0_in_h,
  /* <bf2> */ output mbx5_rq_1_in_h,
  /* <bf1> */ output mbx5_rq_2_in_h,
  /* <be2> */ output mbx5_rq_3_in_h,
  /* <cr1> */  input mcl2_vma_pause_l,
  /* <fk1> */  input mcl6_ebox_cache_l,
  /* <at2> */ output mem_data_to_mem_h,
  /* <ce2> */ output mem_diag_l,
  /* <em2> */  input mem_rd_rq_h,
  /* <dm1> */  input mem_to_c_diag_en_l,
  /* <bv2> */ output mem_to_c_sel_1_h,
  /* <bu2> */ output mem_to_c_sel_2_h,
  /* <fm2> */  input mr_reset_06_h,
  /* <fk2> */  input pag1_pt_cache_l,
  /* <cl1> */  input phase_change_coming_l,
  /* <fl1> */  input pma2_cca_cry_out_l,
  /* <ck1> */  input pma4_pa_34_h,
  /* <cj1> */  input pma4_pa_35_h,
  /* <dp2> */  input pma5_csh_ebox_cyc_l,
  /* <ee1> */  input pma5_csh_writeback_cyc_h,
  /* <fa1> */  input pma5_ebox_paged_l,
  /* <be1> */ output sbus_adr_34_h,
  /* <bd2> */ output sbus_adr_35_h
);

`include "mbx21.svh"

endmodule	// mbx21
