module chx28(
      input  apr_en_refill_ram_wr_h            /* <aj2> */,
      output cam_14_h                          /* <bv2> */,
      output cam_15_h                          /* <bt2> */,
      output cam_16_h                          /* <ck2> */,
      output cam_17_h                          /* <ce2> */,
      output cam_18_h                          /* <cu2> */,
      output cam_19_h                          /* <cs2> */,
      output cam_20_h                          /* <ej1> */,
      output cam_21_h                          /* <ej2> */,
      output cam_22_h                          /* <ff1> */,
      output cam_23_h                          /* <fc1> */,
      output cam_24_h                          /* <fm2> */,
      output cam_25_h                          /* <fk2> */,
      output cam_26_h                          /* <fv2> */,
      output cam_par_h                         /* <fs2> */,
      input  cam_sel_1_h                       /* <cl2> */,
      input  cam_sel_2_h                       /* <bu2> */,
      input  clk_chx_h                         /* <cr2> */,
      output csh_0_00to17_sel_a_l              /* <ap2> */,
      output csh_0_18to35_sel_a_l              /* <cd2> */,
      output csh_0_valid_match_h               /* <cp2> */,
      output csh_0_valid_match_l               /* <cm2> */,
      output csh_0_wd_val_h                    /* <au2> */,
      input  csh_0_wr_en_l                     /* <al1> */,
      output csh_1_00to17_sel_a_l              /* <cv2> */,
      output csh_1_18to35_sel_a_l              /* <ct2> */,
      output csh_1_valid_match_h               /* <cj2> */,
      output csh_1_valid_match_l               /* <bs2> */,
      output csh_1_wd_val_h                    /* <ar2> */,
      input  csh_1_wr_en_l                     /* <am1> */,
      output csh_2_00to17_sel_a_l              /* <en1> */,
      output csh_2_18to35_sel_a_l              /* <ek1> */,
      output csh_2_valid_match_h               /* <fe2> */,
      output csh_2_valid_match_l               /* <ff2> */,
      output csh_2_wd_val_h                    /* <bj2> */,
      input  csh_2_wr_en_l                     /* <aj1> */,
      output csh_3_00to17_sel_a_l              /* <fm1> */,
      output csh_3_18to35_sel_a_l              /* <fj1> */,
      output csh_3_valid_match_h               /* <et2> */,
      output csh_3_valid_match_l               /* <fa1> */,
      output csh_3_wd_val_h                    /* <bh2> */,
      input  csh_3_wr_en_l                     /* <ak2> */,
      output csh_adr_par_bad_l                 /* <fh2> */,
      input  csh_dir_14_0_h                    /* <da1> */,
      input  csh_dir_14_1_h                    /* <cj1> */,
      input  csh_dir_14_2_h                    /* <dl2> */,
      input  csh_dir_14_3_h                    /* <df2> */,
      input  csh_dir_15_0_h                    /* <cm1> */,
      input  csh_dir_15_1_h                    /* <cd1> */,
      input  csh_dir_15_2_h                    /* <dl1> */,
      input  csh_dir_15_3_h                    /* <de1> */,
      input  csh_dir_16_0_h                    /* <cl1> */,
      input  csh_dir_16_1_h                    /* <cc1> */,
      input  csh_dir_16_2_h                    /* <ca1> */,
      input  csh_dir_16_3_h                    /* <dc1> */,
      input  csh_dir_17_0_h                    /* <cp1> */,
      input  csh_dir_17_1_h                    /* <cf1> */,
      input  csh_dir_17_2_h                    /* <ce1> */,
      input  csh_dir_17_3_h                    /* <dd2> */,
      input  csh_dir_18_0_h                    /* <dr1> */,
      input  csh_dir_18_1_h                    /* <dt2> */,
      input  csh_dir_18_2_h                    /* <ef1> */,
      input  csh_dir_18_3_h                    /* <ea1> */,
      input  csh_dir_19_0_h                    /* <dn1> */,
      input  csh_dir_19_1_h                    /* <ds1> */,
      input  csh_dir_19_2_h                    /* <ee2> */,
      input  csh_dir_19_3_h                    /* <ec1> */,
      input  csh_dir_20_0_h                    /* <dj1> */,
      input  csh_dir_20_1_h                    /* <dm1> */,
      input  csh_dir_20_2_h                    /* <du2> */,
      input  csh_dir_20_3_h                    /* <dr2> */,
      input  csh_dir_21_0_h                    /* <dk1> */,
      input  csh_dir_21_1_h                    /* <dm2> */,
      input  csh_dir_21_2_h                    /* <dv2> */,
      input  csh_dir_21_3_h                    /* <ds2> */,
      input  csh_dir_22_0_h                    /* <eh2> */,
      input  csh_dir_22_1_h                    /* <ep2> */,
      input  csh_dir_22_2_h                    /* <fd1> */,
      input  csh_dir_22_3_h                    /* <es2> */,
      input  csh_dir_23_0_h                    /* <ef2> */,
      input  csh_dir_23_1_h                    /* <ep1> */,
      input  csh_dir_23_2_h                    /* <fe1> */,
      input  csh_dir_23_3_h                    /* <er1> */,
      input  csh_dir_24_0_h                    /* <ed1> */,
      input  csh_dir_24_1_h                    /* <ek2> */,
      input  csh_dir_24_2_h                    /* <eu2> */,
      input  csh_dir_24_3_h                    /* <el2> */,
      input  csh_dir_25_0_h                    /* <ee1> */,
      input  csh_dir_25_1_h                    /* <el1> */,
      input  csh_dir_25_2_h                    /* <ev2> */,
      input  csh_dir_25_3_h                    /* <em1> */,
      input  csh_dir_26_0_h                    /* <fd2> */,
      input  csh_dir_26_1_h                    /* <fl2> */,
      input  csh_dir_26_2_h                    /* <fu2> */,
      input  csh_dir_26_3_h                    /* <fk1> */,
      input  csh_dir_par_0_h                   /* <fr2> */,
      input  csh_dir_par_1_h                   /* <fp1> */,
      input  csh_dir_par_2_h                   /* <fn1> */,
      input  csh_dir_par_3_h                   /* <fp2> */,
      output csh_lru_1_h                       /* <br1> */,
      output csh_lru_2_h                       /* <bs1> */,
      input  csh_refill_ram_wr_l               /* <am2> */,
      input  csh_sel_lru_h                     /* <av2> */,
      input  csh_sel_lru_l                     /* <bp2> */,
      input  csh_use_hold_h                    /* <al2> */,
      input  csh_use_wr_en_h                   /* <br2> */,
      input  csh_val_sel_all_h                 /* <ac1> */,
      input  csh_val_wr_data_h                 /* <bk1> */,
      input  csh_val_wr_pulse_l                /* <ak1> */,
      output csh_wd_0_val_h                    /* <bl2> */,
      output csh_wd_1_val_h                    /* <bk2> */,
      output csh_wd_2_val_h                    /* <bf2> */,
      output csh_wd_3_val_h                    /* <bd2> */,
      input  csh_wr_wd_0_en_h                  /* <ae1> */,
      input  csh_wr_wd_1_en_h                  /* <af1> */,
      input  csh_wr_wd_2_en_h                  /* <aa1> */,
      input  csh_wr_wd_3_en_h                  /* <ad1> */,
      input  diag_04_b_h                       /* <ft2> */,
      input  diag_05_b_h                       /* <fs1> */,
      input  diag_06_b_h                       /* <fr1> */,
      input  diag_read_func_17x_l              /* <bn1> */,
      output ebus_d20_e_h                      /* <ch2> */,
      output ebus_d21_e_h                      /* <cf2> */,
      input  force_no_match_h                  /* <fj2> */,
      input  force_valid_match_0_h             /* <cs1> */,
      input  force_valid_match_1_h             /* <ck1> */,
      input  force_valid_match_2_h             /* <dh2> */,
      input  force_valid_match_3_h             /* <dd1> */,
      input  mbx_csh_adr_27_h                  /* <as1> */,
      input  mbx_csh_adr_28_h                  /* <an1> */,
      input  mbx_csh_adr_29_h                  /* <be1> */,
      input  mbx_csh_adr_30_h                  /* <ba1> */,
      input  mbx_csh_adr_31_h                  /* <bp1> */,
      input  mbx_csh_adr_32_h                  /* <bl1> */,
      input  mbx_csh_adr_33_h                  /* <bf1> */,
      input  pma_34_h                          /* <as2> */,
      input  pma_35_h                          /* <be2> */,
      input  pt_14_b_h                         /* <df1> */,
      input  pt_15_b_h                         /* <de2> */,
      input  pt_16_b_h                         /* <cn1> */,
      input  pt_17_b_h                         /* <cr1> */,
      input  pt_18_b_h                         /* <dp2> */,
      input  pt_19_b_h                         /* <dp1> */,
      input  pt_20_b_h                         /* <dj2> */,
      input  pt_21_b_h                         /* <dk2> */,
      input  pt_22_b_h                         /* <es1> */,
      input  pt_23_b_h                         /* <er2> */,
      input  pt_24_b_h                         /* <ed2> */,
      input  pt_25_b_h                         /* <em2> */,
      input  pt_26_b_h                         /* <fl1> */,
      input  vma_18_a_h                        /* <af2> */,
      input  vma_19_a_h                        /* <ae2> */,
      input  vma_20_a_h                        /* <ad2> */,
      input  vma_27_g_h                        /* <ar1> */,
      input  vma_28_g_h                        /* <ap1> */,
      input  vma_29_g_h                        /* <bd1> */,
      input  vma_30_g_h                        /* <bc1> */,
      input  vma_31_g_h                        /* <bm2> */,
      input  vma_32_g_h                        /* <bm1> */,
      input  vma_33_g_h                        /* <bj1> */
);

`include "chx28nets.svh"

endmodule	// chx28
