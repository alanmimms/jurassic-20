`ifndef __LOGIC_SVH__
`define __LOGIC_SVH__ 1

// MC10141 mode
typedef enum bit [1:0] {LOAD, SHIFTL, SHIFTR, HOLD} tMode141;

`endif
