module just_a_wire(input bit b, output bit q);
  assign q = b;
endmodule // just_a_wire
