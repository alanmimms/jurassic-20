module con;
`include "con.svh"
endmodule	// con
