module apr34(
      output apr2_c_dir_p_err_h                /* <ep1> */,
      output apr2_clk_c_h                      /* <dj2> */,
      output apr2_wr_bad_adr_par_l             /* <ch2> */,
      output apr3_coni_or_datai_l              /* <bj2> */,
      output apr3_cono_or_datao_h              /* <bm1> */,
      output apr3_fetch_comp_h                 /* <br2> */,
      output apr3_fm_extended_h                /* <ce2> */,
      output apr3_fm_odd_parity_h              /* <dd1> */,
      output apr3_read_comp_h                  /* <cj2> */,
      input  apr3_spare_l                      /* <df1> */,
      output apr3_user_comp_h                  /* <ce1> */,
      output apr3_write_comp_h                 /* <ck1> */,
      output apr4_ac_09_l                      /* <ef1> */,
      output apr4_ac_10_l                      /* <ba1> */,
      output apr4_ac_11_l                      /* <fd1> */,
      output apr4_ac_12_l                      /* <ft2> */,
      output apr5_mbox_ctl_06_l                /* <al1> */,
      output apr5_pt_dir_wr_l                  /* <bd2> */,
      output apr5_pt_wr_l                      /* <bc1> */,
      output apr5_set_page_fail_l              /* <bd1> */,
      output apr5_wr_pt_sel_0_h                /* <bj1> */,
      output apr5_wr_pt_sel_1_h                /* <bf1> */,
      output apr5_wr_pt_sel_1_l                /* <al2> */,
      output apr6_ebox_cca_h                   /* <cc1> */,
      output apr6_ebox_cca_l                   /* <ac1> */,
      output apr6_ebox_ebr_h                   /* <cd1> */,
      output apr6_ebox_era_l                   /* <ad1> */,
      output apr6_ebox_load_reg_l              /* <dd2> */,
      output apr6_ebox_read_reg_h              /* <ap2> */,
      output apr6_ebox_read_reg_l              /* <dc1> */,
      output apr6_ebox_sbus_diag_h             /* <cu2> */,
      output apr6_ebox_ubr_h                   /* <cd2> */,
      output apr_any_ebox_err_flg_h            /* <cj1> */,
      output apr_apr_interrupt_l               /* <cl1> */,
      output apr_ebox_disable_cs_h             /* <cf1> */,
      output apr_ebox_era_h                    /* <au2> */,
      output apr_ebox_sbus_diag_l              /* <cn1> */,
      output apr_ebox_send_f02_h               /* <bu2> */,
      output apr_ebox_spare_h                  /* <as2> */,
      output apr_ebus_demand_h                 /* <bp1> */,
      output apr_ebus_f01_e_h                  /* <bv2> */,
      output apr_ebus_req_l                    /* <be2> */,
      output apr_ebus_return_h                 /* <bp2> */,
      output apr_en_refill_ram_wr_h            /* <at2> */,
      output apr_fm_36_h                       /* <de2> */,
      output apr_fm_adr_10_h                   /* <bt2> */,
      output apr_fm_adr_1_h                    /* <cv2> */,
      output apr_fm_adr_2_h                    /* <av2> */,
      output apr_fm_adr_4_h                    /* <ca1> */,
      output apr_fm_block_1_h                  /* <cf2> */,
      output apr_fm_block_2_h                  /* <br1> */,
      output apr_fm_block_4_h                  /* <be1> */,
      output apr_mb_par_err_l                  /* <fa1> */,
      output apr_mbox_ctl_03_h                 /* <bh2> */,
      output apr_mbox_ctl_06_h                 /* <bf2> */,
      output apr_nxm_err_l                     /* <bs1> */,
      output apr_s_adr_p_err_l                 /* <ae2> */,
      output apr_sbus_err_l                    /* <bs2> */,
      input  clk3_apr_h                        /* <cr2> */,
      input  con_condSlebus_ctl_l              /* <bk1> */,
      input  con_condSlmbox_ctl_l              /* <af1> */,
      input  con_datao_apr_l                   /* <dk2> */,
      input  con_fm_write_par_l                /* <ck2> */,
      input  con_load_ac_blocks_l              /* <er2> */,
      input  con_sel_clr_h                     /* <dt2> */,
      input  con_sel_dis_h                     /* <ej2> */,
      input  con_sel_en_l                      /* <ek2> */,
      input  con_sel_set_l                     /* <du2> */,
      input  con_wr_even_par_adr_h             /* <ad2> */,
      input  cram_Nr_00_d_h                    /* <aa1> */,
      input  cram_Nr_01_d_h                    /* <an1> */,
      input  cram_Nr_02_d_h                    /* <ep2> */,
      input  cram_Nr_03_d_h                    /* <ap1> */,
      input  cram_Nr_04_d_h                    /* <ar2> */,
      input  cram_Nr_05_d_h                    /* <as1> */,
      input  cram_Nr_06_d_h                    /* <aj1> */,
      input  cram_Nr_07_d_h                    /* <ak2> */,
      input  cram_Nr_08_d_h                    /* <am1> */,
      input  cram_adb_sel_1_h                  /* <fs2> */,
      input  cram_adb_sel_2_h                  /* <fr2> */,
      input  cram_fm_adr_sel_1_h               /* <ef2> */,
      input  cram_fm_adr_sel_2s_h              /* <ee1> */,
      input  cram_fm_adr_sel_4_h               /* <ed2> */,
      input  ctl3_diag_rd_func_11x_l           /* <bn1> */,
      input  diag_04_b_h                       /* <bl2> */,
      input  diag_05_b_h                       /* <bm2> */,
      input  diag_06_b_h                       /* <bl1> */,
      output ebus_d01_e_h                      /* <cm1> */,
      output ebus_d06_e_h                      /* <cm2> */,
      output ebus_d07_e_h                      /* <cp1> */,
      output ebus_d08_e_h                      /* <cp2> */,
      output ebus_d09_e_h                      /* <cl2> */,
      output ebus_d10_e_h                      /* <cr1> */,
      output ebus_d11_e_h                      /* <ds1> */,
      output ebus_d12_e_h                      /* <cs1> */,
      output ebus_d13_e_h                      /* <cs2> */,
      output ebus_d14_e_h                      /* <dk1> */,
      output ebus_d15_e_h                      /* <dl1> */,
      output ebus_d16_e_h                      /* <dl2> */,
      output ebus_d17_e_h                      /* <dp1> */,
      input  edp_fm_parity_00to05_h            /* <fl2> */,
      input  edp_fm_parity_06to11_h            /* <fk2> */,
      input  edp_fm_parity_12to17_h            /* <fj2> */,
      input  edp_fm_parity_18to23_h            /* <ff2> */,
      input  edp_fm_parity_24to29_h            /* <ff1> */,
      input  edp_fm_parity_30to35_h            /* <fe2> */,
      input  ir_ac_09_h                        /* <ed1> */,
      input  ir_ac_10_h                        /* <ec1> */,
      input  ir_ac_11_h                        /* <ea1> */,
      input  ir_ac_12_h                        /* <dv2> */,
      input  mbox_adr_par_err_l                /* <ae1> */,
      input  mbox_mb_par_err_l                 /* <fc1> */,
      input  mbox_nxm_err_l                    /* <el2> */,
      input  mbox_sbus_err_l                   /* <el1> */,
      input  mbx1_cca_req_l                    /* <em2> */,
      input  mbx5_csh_adr_par_err_l            /* <dr2> */,
      input  mcl1_memSlreg_func_l              /* <aj2> */,
      input  mcl1_req_en_l                     /* <ak1> */,
      input  mcl4_load_vma_context_l           /* <af2> */,
      input  mcl4_vma_prev_en_h                /* <am2> */,
      input  mcl4_xr_previous_h                /* <fm1> */,
      input  mcl6_ebox_map_h                   /* <ar1> */,
      input  mr_reset_02_h                     /* <ah2> */,
      input  pi3_apr_pia_01_h                  /* <da1> */,
      input  pi3_apr_pia_02_h                  /* <dh2> */,
      input  pi3_apr_pia_04_h                  /* <ct2> */,
      input  pwr_warn_e_h                      /* <en1> */,
      input  shm1_ar_extended_h                /* <er1> */,
      input  shm1_ar_par_odd_b_h               /* <eu2> */,
      input  shm1_xr_01_h                      /* <fu2> */,
      input  shm1_xr_02_h                      /* <fp2> */,
      input  shm1_xr_04_h                      /* <et2> */,
      input  shm1_xr_10_h                      /* <ej1> */,
      input  vma1_vma_32_b_h                   /* <eh2> */,
      input  vma1_vma_33_b_h                   /* <es1> */,
      input  vma1_vma_34_b_h                   /* <fp1> */,
      input  vma1_vma_35_b_h                   /* <fv2> */
);

`include "apr34nets.svh"

endmodule	// apr34
