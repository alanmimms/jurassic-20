module delay_line(input bit in, output bit out);
  assign out = in;
endmodule // delay_line
