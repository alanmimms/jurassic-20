module mb014(
      input  ar_12_a_h                         /* <fc1> */,
      input  ar_13_a_h                         /* <fd1> */,
      input  ar_14_a_h                         /* <eu2> */,
      input  ar_15_a_h                         /* <ev2> */,
      input  ar_16_a_h                         /* <cv2> */,
      input  ar_17_a_h                         /* <bu2> */,
      input  ar_30_a_h                         /* <dd2> */,
      input  ar_31_a_h                         /* <cs2> */,
      input  ar_32_a_h                         /* <bp1> */,
      input  ar_33_a_h                         /* <bj2> */,
      input  ar_34_a_h                         /* <bm2> */,
      input  ar_35_a_h                         /* <bf1> */,
      input  cache_data_12_a_h                 /* <er2> */,
      input  cache_data_13_a_h                 /* <ef1> */,
      input  cache_data_14_a_h                 /* <ff2> */,
      input  cache_data_15_a_h                 /* <er1> */,
      input  cache_data_16_a_h                 /* <cr1> */,
      input  cache_data_17_a_h                 /* <cm2> */,
      input  cache_data_30_a_h                 /* <dk2> */,
      input  cache_data_31_a_h                 /* <dk1> */,
      input  cache_data_32_a_h                 /* <am1> */,
      input  cache_data_33_a_h                 /* <ak1> */,
      input  cache_data_34_a_h                 /* <ar1> */,
      input  cache_data_35_a_h                 /* <ap1> */,
      input  cbus_d12_re_h                     /* <cj1> */,
      output cbus_d12_te_h                     /* <ee1> */,
      input  cbus_d13_re_h                     /* <cj2> */,
      output cbus_d13_te_h                     /* <ee2> */,
      input  cbus_d14_re_h                     /* <bs2> */,
      output cbus_d14_te_h                     /* <el2> */,
      input  cbus_d15_re_h                     /* <bc1> */,
      output cbus_d15_te_h                     /* <em1> */,
      input  cbus_d16_re_h                     /* <br1> */,
      output cbus_d16_te_h                     /* <df1> */,
      input  cbus_d17_re_h                     /* <bd2> */,
      output cbus_d17_te_h                     /* <dl2> */,
      input  cbus_d30_re_h                     /* <ch2> */,
      output cbus_d30_te_h                     /* <dn1> */,
      input  cbus_d31_re_h                     /* <cf1> */,
      output cbus_d31_te_h                     /* <dm2> */,
      input  cbus_d32_re_h                     /* <be2> */,
      output cbus_d32_te_h                     /* <ah2> */,
      input  cbus_d33_re_h                     /* <bj1> */,
      output cbus_d33_te_h                     /* <af2> */,
      input  cbus_d34_re_h                     /* <be1> */,
      output cbus_d34_te_h                     /* <aj2> */,
      input  cbus_d35_re_h                     /* <bl1> */,
      output cbus_d35_te_h                     /* <ak2> */,
      input  ccl_ccw_buf_wr_l                  /* <fk1> */,
      input  ccl_ch_buf_en_l                   /* <ae2> */,
      input  ccl_mix_mb_sel_h                  /* <es1> */,
      input  ccw_buf_12_in_h                   /* <fl1> */,
      input  ccw_buf_13_in_h                   /* <fm2> */,
      input  ccw_buf_14_in_h                   /* <fh2> */,
      input  ccw_buf_15_in_h                   /* <fj2> */,
      input  ccw_buf_16_in_h                   /* <cl2> */,
      input  ccw_buf_17_in_h                   /* <cl1> */,
      input  ccw_buf_30_in_h                   /* <ck2> */,
      input  ccw_buf_31_in_h                   /* <ck1> */,
      input  ccw_buf_32_in_h                   /* <at2> */,
      input  ccw_buf_33_in_h                   /* <as1> */,
      input  ccw_buf_34_in_h                   /* <ap2> */,
      input  ccw_buf_35_in_h                   /* <am2> */,
      input  ccw_buf_adr_0_h                   /* <fk2> */,
      input  ccw_buf_adr_1_h                   /* <fj1> */,
      input  ccw_buf_adr_2_h                   /* <fl2> */,
      input  ccw_buf_adr_3_h                   /* <fm1> */,
      output ccw_mix_12_h                      /* <ek2> */,
      output ccw_mix_13_h                      /* <eh2> */,
      output ccw_mix_14_h                      /* <ff1> */,
      output ccw_mix_15_h                      /* <es2> */,
      output ccw_mix_16_h                      /* <cp2> */,
      output ccw_mix_17_h                      /* <cn1> */,
      output ccw_mix_30_h                      /* <dl1> */,
      output ccw_mix_31_h                      /* <dh2> */,
      output ccw_mix_32_h                      /* <al2> */,
      output ccw_mix_33_h                      /* <al1> */,
      output ccw_mix_34_h                      /* <as2> */,
      output ccw_mix_35_h                      /* <ar2> */,
      input  ch_buf_wr_05_l                    /* <aj1> */,
      input  ch_buf_wr_2_l                     /* <ep1> */,
      input  ch_reverse_h                      /* <bd1> */,
      input  ch_t0_l                           /* <fs2> */,
      input  ch_t2_l                           /* <af1> */,
      input  clk_mb_12_h                       /* <cr2> */,
      input  con_ki10_paging_mode_l            /* <ek1> */,
      input  crc_buf_mb_sel_h                  /* <dt2> */,
      input  crc_cbus_out_hold_h               /* <fu2> */,
      input  crc_ch_buf_adr_0_h                /* <fp2> */,
      input  crc_ch_buf_adr_1_h                /* <fr2> */,
      input  crc_ch_buf_adr_2_h                /* <fp1> */,
      input  crc_ch_buf_adr_3_h                /* <de1> */,
      input  crc_ch_buf_adr_4_h                /* <dj1> */,
      input  crc_ch_buf_adr_5_h                /* <de2> */,
      input  crc_ch_buf_adr_6_h                /* <ae1> */,
      input  mb0_hold_in_h                     /* <ad2> */,
      input  mb1_hold_in_h                     /* <ad1> */,
      input  mb2_hold_in_h                     /* <aa1> */,
      input  mb3_hold_in_h                     /* <ac1> */,
      output mb_12_h                           /* <fd2> */,
      output mb_12to17_par_odd_h               /* <ds2> */,
      output mb_13_h                           /* <dr2> */,
      output mb_14_h                           /* <dp2> */,
      output mb_15_h                           /* <dm1> */,
      output mb_16_h                           /* <dr1> */,
      output mb_17_h                           /* <dp1> */,
      output mb_30_h                           /* <av2> */,
      output mb_30to35_par_odd_h               /* <au2> */,
      output mb_31_h                           /* <ba1> */,
      output mb_32_h                           /* <cd2> */,
      output mb_33_h                           /* <cd1> */,
      output mb_34_h                           /* <ca1> */,
      output mb_35_h                           /* <bv2> */,
      input  mb_in_sel_1_h                     /* <ej1> */,
      input  mb_in_sel_2_h                     /* <el1> */,
      input  mb_in_sel_4_h                     /* <ep2> */,
      input  mb_sel_1_en_h                     /* <fr1> */,
      input  mb_sel_2_en_h                     /* <ft2> */,
      input  mb_sel_hold_h                     /* <fv2> */,
      input  mem_data_in_12_h                  /* <em2> */,
      input  mem_data_in_13_h                  /* <ej2> */,
      input  mem_data_in_14_h                  /* <ea1> */,
      input  mem_data_in_15_h                  /* <dv2> */,
      input  mem_data_in_16_h                  /* <cp1> */,
      input  mem_data_in_17_h                  /* <cm1> */,
      input  mem_data_in_30_h                  /* <dj2> */,
      input  mem_data_in_31_h                  /* <df2> */,
      input  mem_data_in_32_h                  /* <bm1> */,
      input  mem_data_in_33_h                  /* <bk2> */,
      input  mem_data_in_34_h                  /* <bl2> */,
      input  mem_data_in_35_h                  /* <bk1> */,
      input  mem_to_c_en_l                     /* <ed2> */,
      input  mem_to_c_sel_1_h                  /* <ed1> */,
      input  mem_to_c_sel_2_h                  /* <ds1> */,
      output mem_to_cache_12_h                 /* <en1> */,
      output mem_to_cache_13_h                 /* <ef2> */,
      output mem_to_cache_14_h                 /* <ec1> */,
      output mem_to_cache_15_h                 /* <du2> */,
      output mem_to_cache_16_h                 /* <cf2> */,
      output mem_to_cache_17_h                 /* <cc1> */,
      output mem_to_cache_30_h                 /* <cs1> */,
      output mem_to_cache_31_h                 /* <dd1> */,
      output mem_to_cache_32_h                 /* <br2> */,
      output mem_to_cache_33_h                 /* <bf2> */,
      output mem_to_cache_34_h                 /* <bp2> */,
      output mem_to_cache_35_h                 /* <bh2> */,
      input  nxm_any_l                         /* <fs1> */,
      output pt_in_12_h                        /* <fe1> */,
      output pt_in_13_h                        /* <fe2> */,
      output pt_in_14_h                        /* <fa1> */,
      output pt_in_15_h                        /* <et2> */,
      output pt_in_16_h                        /* <dc1> */,
      output pt_in_17_h                        /* <da1> */,
      output pt_in_30_h                        /* <cu2> */,
      output pt_in_31_h                        /* <ct2> */,
      output pt_in_32_h                        /* <ce1> */,
      output pt_in_33_h                        /* <ce2> */,
      output pt_in_34_h                        /* <bs1> */,
      output pt_in_35_h                        /* <bt2> */
);

`include "mb014nets.svh"

endmodule	// mb014
