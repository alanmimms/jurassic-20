module vma;
`include "vma.svh"
endmodule	// vma
