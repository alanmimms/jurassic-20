module clk32(
  /* <eh2> */  input apr3_fm_odd_parity_h,
  /* <dm1> */  input apr5_pt_dir_wr_l,
  /* <dj2> */  input apr5_pt_wr_l,
  /* <ea1> */  input apr5_set_page_fail_l,
  /* <cp2> */  input apr_apr_par_chk_en_l,
  /* <dd2> */ output clk1_chc_h,
  /* <cr2> */  input clk1_clk_h,
  /* <fr2> */ output clk1_clk_out_h,
  /* <fd2> */ output clk1_csh_h,
  /* <es2> */ output clk1_mbc_h,
  /* <ef2> */ output clk1_mbox_13_a_h,
  /* <ee2> */ output clk1_mbox_14_a_h,
  /* <er2> */ output clk1_mbx_h,
  /* <fs2> */ output clk1_mtr_h,
  /* <ff2> */ output clk1_pma_h,
  /* <dn1> */ output clk2_pt_dir_wr_l,
  /* <dl2> */ output clk2_pt_wr_l,
  /* <cs2> */ output clk3_apr_h,
  /* <am1> */ output clk3_arSlarx_mem_load_h,
  /* <ba1> */ output clk3_ebox_sync_b_l,
  /* <bc1> */ output clk3_ebox_sync_c_l,
  /* <au2> */ output clk3_ebox_sync_d_l,
  /* <em1> */  input clk3_fs_en_a_h,
  /* <el1> */  input clk3_fs_en_b_h,
  /* <el2> */  input clk3_fs_en_c_h,
  /* <ek1> */  input clk3_fs_en_d_h,
  /* <ej1> */  input clk3_fs_en_e_l,
  /* <ej2> */  input clk3_fs_en_f_l,
  /* <ek2> */  input clk3_fs_en_g_l,
  /* <cf2> */ output clk3_mcl_h,
  /* <cd2> */ output clk3_scd_h,
  /* <cj2> */ output clk3_vma_h,
  /* <dm2> */ output clk4_ebox_cyc_abort_h,
  /* <bm1> */ output clk4_ebox_req_h,
  /* <aj1> */ output clk4_ebox_req_l,
  /* <bm2> */ output clk4_force_1777_h,
  /* <cf1> */ output clk4_pf_disp_07_h,
  /* <cc1> */ output clk4_pf_disp_08_h,
  /* <cm1> */ output clk4_pf_disp_09_h,
  /* <ch2> */ output clk4_pf_disp_10_h,
  /* <am2> */ output clk4_resp_mbox_h,
  /* <fj2> */ output clk_10_11_clk_h,
  /* <df2> */ output clk_ccl_h,
  /* <dp2> */ output clk_ccw_h,
  /* <fe2> */ output clk_chx_h,
  /* <ck2> */ output clk_con_h,
  /* <ap2> */ output clk_cra_h,
  /* <de2> */ output clk_crc_h,
  /* <as2> */ output clk_crm_00_h,
  /* <ar2> */ output clk_crm_04_h,
  /* <af2> */ output clk_crm_08_h,
  /* <ae2> */ output clk_crm_12_h,
  /* <ad2> */ output clk_crm_16_h,
  /* <av2> */ output clk_ebox_sync_a_l,
  /* <bk1> */ output clk_ebus_clk_h,
  /* <dt2> */ output clk_ebus_reset_e_h,
  /* <bd2> */ output clk_edp_00_h,
  /* <be2> */ output clk_edp_06_h,
  /* <bf2> */ output clk_edp_12_h,
  /* <bp2> */ output clk_edp_18_h,
  /* <br2> */ output clk_edp_24_h,
  /* <bs2> */ output clk_edp_30_h,
  /* <bj1> */ output clk_error_stop_h,
  /* <ak2> */ output clk_instr_1777_l,
  /* <ce2> */ output clk_ir_h,
  /* <ed2> */ output clk_mb_00_h,
  /* <ds2> */ output clk_mb_06_h,
  /* <dr2> */ output clk_mb_12_h,
  /* <bl1> */ output clk_mb_xfer_h,
  /* <al1> */ output clk_mb_xfer_l,
  /* <ep2> */ output clk_mbz_h,
  /* <an1> */ output clk_page_error_h,
  /* <fp2> */ output clk_pi_h,
  /* <at2> */ output clk_sbr_call_h,
  /* <ca1> */ output clk_sbus_clk_h,
  /* <bl2> */  input con_ar_from_ebus_h,
  /* <cr1> */  input con_ar_loaded_l,
  /* <cp1> */  input con_arx_loaded_l,
  /* <dh2> */  input con_cono_200000_h,
  /* <cu2> */  input con_delay_req_h,
  /* <fk1> */  input con_load_dram_h,
  /* <cn1> */  input con_mbox_wait_l,
  /* <fn1> */  input cram_mem_02_a_h,
  /* <fl1> */  input cram_par_16_h,
  /* <da1> */  input cram_t_00_h,
  /* <cv2> */  input cram_t_01_h,
  /* <fh2> */  input crobar_e_h,
  /* <ac1> */  input csh2_ebox_retry_req_l,
  /* <ak1> */  input csh2_mbox_resp_in_h,
  /* <bk2> */  input csh4_ebox_t0_in_h,
  /* <aj2> */  input csh6_page_fail_hold_h,
  /* <bj2> */  input ctl3_diag_clk_edp_h,
  /* <fk2> */  input ctl3_diag_ctl_func_00x_l,
  /* <fm1> */  input ctl3_diag_ld_func_04x_l,
  /* <ec1> */  input deskew_clk_h,
  /* <du2> */  input diag_channel_clk_stop_h,
  /* <bn1> */  input diag_read_func_10x_l,
  /* <fj1> */  input dram_odd_parity_h,
  /* <cl1> */ output ebus_d30_e_h,
  /* <cl2> */ output ebus_d31_e_h,
  /* <dc1> */ output ebus_d32_e_h,
  /* <dj1> */ output ebus_d33_e_h,
  /* <dk1> */ output ebus_d34_e_h,
  /* <dl1> */ output ebus_d35_e_h,
  /* <bu2> */  input ebus_ds04_e_h,
  /* <bv2> */  input ebus_ds05_e_h,
  /* <bt2> */  input ebus_ds06_e_h,
  /* <fv2> */  input external_clk_h,
  /* <aa1> */  input mcl5_mbox_cyc_req_l,
  /* <fc1> */ output mr_reset_01_h,
  /* <fa1> */ output mr_reset_02_h,
  /* <et2> */ output mr_reset_04_h,
  /* <eu2> */ output mr_reset_05_h,
  /* <em2> */ output mr_reset_06_h,
  /* <en1> */  input pag4_pf_ebox_handle_h,
  /* <ct2> */  input shm1_ar_par_odd_h,
  /* <cm2> */  input shm1_arx_par_odd_h,
  /* <fm2> */  input synchronize_clk_h,
  /* <al2> */  input vma1_ac_ref_h
);

`include "clk32.svh"

endmodule	// clk32
