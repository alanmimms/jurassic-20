module chx28(
  /* <aj2> */  input apr_en_refill_ram_wr_h,
  /* <bv2> */ output cam_14_h,
  /* <bt2> */ output cam_15_h,
  /* <ck2> */ output cam_16_h,
  /* <ce2> */ output cam_17_h,
  /* <cu2> */ output cam_18_h,
  /* <cs2> */ output cam_19_h,
  /* <ej1> */ output cam_20_h,
  /* <ej2> */ output cam_21_h,
  /* <ff1> */ output cam_22_h,
  /* <fc1> */ output cam_23_h,
  /* <fm2> */ output cam_24_h,
  /* <fk2> */ output cam_25_h,
  /* <fv2> */ output cam_26_h,
  /* <fs2> */ output cam_par_h,
  /* <cl2> */  input cam_sel_1_h,
  /* <bu2> */  input cam_sel_2_h,
  /* <cr2> */  input clk_chx_h,
  /* <ap2> */ output csh_0_00to17_sel_a_l,
  /* <cd2> */ output csh_0_18to35_sel_a_l,
  /* <cp2> */ output csh_0_valid_match_h,
  /* <cm2> */ output csh_0_valid_match_l,
  /* <au2> */ output csh_0_wd_val_h,
  /* <al1> */  input csh_0_wr_en_l,
  /* <cv2> */ output csh_1_00to17_sel_a_l,
  /* <ct2> */ output csh_1_18to35_sel_a_l,
  /* <cj2> */ output csh_1_valid_match_h,
  /* <bs2> */ output csh_1_valid_match_l,
  /* <ar2> */ output csh_1_wd_val_h,
  /* <am1> */  input csh_1_wr_en_l,
  /* <en1> */ output csh_2_00to17_sel_a_l,
  /* <ek1> */ output csh_2_18to35_sel_a_l,
  /* <fe2> */ output csh_2_valid_match_h,
  /* <ff2> */ output csh_2_valid_match_l,
  /* <bj2> */ output csh_2_wd_val_h,
  /* <aj1> */  input csh_2_wr_en_l,
  /* <fm1> */ output csh_3_00to17_sel_a_l,
  /* <fj1> */ output csh_3_18to35_sel_a_l,
  /* <et2> */ output csh_3_valid_match_h,
  /* <fa1> */ output csh_3_valid_match_l,
  /* <bh2> */ output csh_3_wd_val_h,
  /* <ak2> */  input csh_3_wr_en_l,
  /* <fh2> */ output csh_adr_par_bad_l,
  /* <da1> */  input csh_dir_14_0_h,
  /* <cj1> */  input csh_dir_14_1_h,
  /* <dl2> */  input csh_dir_14_2_h,
  /* <df2> */  input csh_dir_14_3_h,
  /* <cm1> */  input csh_dir_15_0_h,
  /* <cd1> */  input csh_dir_15_1_h,
  /* <dl1> */  input csh_dir_15_2_h,
  /* <de1> */  input csh_dir_15_3_h,
  /* <cl1> */  input csh_dir_16_0_h,
  /* <cc1> */  input csh_dir_16_1_h,
  /* <ca1> */  input csh_dir_16_2_h,
  /* <dc1> */  input csh_dir_16_3_h,
  /* <cp1> */  input csh_dir_17_0_h,
  /* <cf1> */  input csh_dir_17_1_h,
  /* <ce1> */  input csh_dir_17_2_h,
  /* <dd2> */  input csh_dir_17_3_h,
  /* <dr1> */  input csh_dir_18_0_h,
  /* <dt2> */  input csh_dir_18_1_h,
  /* <ef1> */  input csh_dir_18_2_h,
  /* <ea1> */  input csh_dir_18_3_h,
  /* <dn1> */  input csh_dir_19_0_h,
  /* <ds1> */  input csh_dir_19_1_h,
  /* <ee2> */  input csh_dir_19_2_h,
  /* <ec1> */  input csh_dir_19_3_h,
  /* <dj1> */  input csh_dir_20_0_h,
  /* <dm1> */  input csh_dir_20_1_h,
  /* <du2> */  input csh_dir_20_2_h,
  /* <dr2> */  input csh_dir_20_3_h,
  /* <dk1> */  input csh_dir_21_0_h,
  /* <dm2> */  input csh_dir_21_1_h,
  /* <dv2> */  input csh_dir_21_2_h,
  /* <ds2> */  input csh_dir_21_3_h,
  /* <eh2> */  input csh_dir_22_0_h,
  /* <ep2> */  input csh_dir_22_1_h,
  /* <fd1> */  input csh_dir_22_2_h,
  /* <es2> */  input csh_dir_22_3_h,
  /* <ef2> */  input csh_dir_23_0_h,
  /* <ep1> */  input csh_dir_23_1_h,
  /* <fe1> */  input csh_dir_23_2_h,
  /* <er1> */  input csh_dir_23_3_h,
  /* <ed1> */  input csh_dir_24_0_h,
  /* <ek2> */  input csh_dir_24_1_h,
  /* <eu2> */  input csh_dir_24_2_h,
  /* <el2> */  input csh_dir_24_3_h,
  /* <ee1> */  input csh_dir_25_0_h,
  /* <el1> */  input csh_dir_25_1_h,
  /* <ev2> */  input csh_dir_25_2_h,
  /* <em1> */  input csh_dir_25_3_h,
  /* <fd2> */  input csh_dir_26_0_h,
  /* <fl2> */  input csh_dir_26_1_h,
  /* <fu2> */  input csh_dir_26_2_h,
  /* <fk1> */  input csh_dir_26_3_h,
  /* <fr2> */  input csh_dir_par_0_h,
  /* <fp1> */  input csh_dir_par_1_h,
  /* <fn1> */  input csh_dir_par_2_h,
  /* <fp2> */  input csh_dir_par_3_h,
  /* <br1> */ output csh_lru_1_h,
  /* <bs1> */ output csh_lru_2_h,
  /* <am2> */  input csh_refill_ram_wr_l,
  /* <av2> */  input csh_sel_lru_h,
  /* <bp2> */  input csh_sel_lru_l,
  /* <al2> */  input csh_use_hold_h,
  /* <br2> */  input csh_use_wr_en_h,
  /* <ac1> */  input csh_val_sel_all_h,
  /* <bk1> */  input csh_val_wr_data_h,
  /* <ak1> */  input csh_val_wr_pulse_l,
  /* <bl2> */ output csh_wd_0_val_h,
  /* <bk2> */ output csh_wd_1_val_h,
  /* <bf2> */ output csh_wd_2_val_h,
  /* <bd2> */ output csh_wd_3_val_h,
  /* <ae1> */  input csh_wr_wd_0_en_h,
  /* <af1> */  input csh_wr_wd_1_en_h,
  /* <aa1> */  input csh_wr_wd_2_en_h,
  /* <ad1> */  input csh_wr_wd_3_en_h,
  /* <bn1> */  input diag_read_func_17x_l,
  /* <ch2> */ output ebus_d20_e_h,
  /* <cf2> */ output ebus_d21_e_h,
  /* <fj2> */  input force_no_match_h,
  /* <cs1> */  input force_valid_match_0_h,
  /* <ck1> */  input force_valid_match_1_h,
  /* <dh2> */  input force_valid_match_2_h,
  /* <dd1> */  input force_valid_match_3_h,
  /* <as1> */  input mbx_csh_adr_27_h,
  /* <an1> */  input mbx_csh_adr_28_h,
  /* <be1> */  input mbx_csh_adr_29_h,
  /* <ba1> */  input mbx_csh_adr_30_h,
  /* <bp1> */  input mbx_csh_adr_31_h,
  /* <bl1> */  input mbx_csh_adr_32_h,
  /* <bf1> */  input mbx_csh_adr_33_h,
  /* <as2> */  input pma_34_h,
  /* <be2> */  input pma_35_h,
  /* <df1> */  input pt_14_b_h,
  /* <de2> */  input pt_15_b_h,
  /* <cn1> */  input pt_16_b_h,
  /* <cr1> */  input pt_17_b_h,
  /* <dp2> */  input pt_18_b_h,
  /* <dp1> */  input pt_19_b_h,
  /* <dj2> */  input pt_20_b_h,
  /* <dk2> */  input pt_21_b_h,
  /* <es1> */  input pt_22_b_h,
  /* <er2> */  input pt_23_b_h,
  /* <ed2> */  input pt_24_b_h,
  /* <em2> */  input pt_25_b_h,
  /* <fl1> */  input pt_26_b_h,
  /* <af2> */  input vma_18_a_h,
  /* <ae2> */  input vma_19_a_h,
  /* <ad2> */  input vma_20_a_h,
  /* <ar1> */  input vma_27_g_h,
  /* <ap1> */  input vma_28_g_h,
  /* <bd1> */  input vma_29_g_h,
  /* <bc1> */  input vma_30_g_h,
  /* <bm2> */  input vma_31_g_h,
  /* <bm1> */  input vma_32_g_h,
  /* <bj1> */  input vma_33_g_h
);

`include "chx28nets.svh"

endmodule	// chx28
