module ird;
`include "ird.svh"
endmodule	// ird
