module shm46(
  /* <ej2> */  input ar_00_b_h,
  /* <em1> */  input ar_01_b_h,
  /* <es1> */  input ar_02_b_h,
  /* <er2> */  input ar_03_b_h,
  /* <ek2> */  input ar_04_b_h,
  /* <ep1> */  input ar_05_b_h,
  /* <ev2> */  input ar_06_b_h,
  /* <fr2> */  input ar_07_b_h,
  /* <ep2> */  input ar_08_b_h,
  /* <em2> */  input ar_09_b_h,
  /* <ff2> */  input ar_10_b_h,
  /* <fu2> */  input ar_11_b_h,
  /* <ej1> */  input ar_12_b_h,
  /* <ee1> */  input ar_13_b_h,
  /* <fk1> */  input ar_14_b_h,
  /* <fj1> */  input ar_15_b_h,
  /* <ef2> */  input ar_16_b_h,
  /* <dp2> */  input ar_17_b_h,
  /* <es2> */  input ar_18_b_h,
  /* <fp2> */  input ar_19_b_h,
  /* <ee2> */  input ar_20_b_h,
  /* <er1> */  input ar_21_b_h,
  /* <fm2> */  input ar_22_b_h,
  /* <fs1> */  input ar_23_b_h,
  /* <fj2> */  input ar_24_b_h,
  /* <el2> */  input ar_25_b_h,
  /* <fr1> */  input ar_26_b_h,
  /* <fs2> */  input ar_27_b_h,
  /* <fk2> */  input ar_28_b_h,
  /* <fl2> */  input ar_29_b_h,
  /* <fp1> */  input ar_30_b_h,
  /* <fv2> */  input ar_31_b_h,
  /* <el1> */  input ar_32_b_h,
  /* <eu2> */  input ar_33_b_h,
  /* <fm1> */  input ar_34_b_h,
  /* <fd1> */  input ar_35_b_h,
  /* <du2> */  input arx_00_a_h,
  /* <dm2> */  input arx_01_a_h,
  /* <cr1> */  input arx_02_h,
  /* <cm2> */  input arx_03_h,
  /* <dl1> */  input arx_04_h,
  /* <cl1> */  input arx_05_h,
  /* <cj2> */  input arx_06_a_h,
  /* <cj1> */  input arx_07_a_h,
  /* <ce1> */  input arx_08_h,
  /* <ce2> */  input arx_09_h,
  /* <cd2> */  input arx_10_h,
  /* <df2> */  input arx_11_h,
  /* <ek1> */  input arx_12_a_h,
  /* <eh2> */  input arx_13_a_h,
  /* <dv2> */  input arx_14_h,
  /* <ff1> */  input arx_15_h,
  /* <ds2> */  input arx_16_h,
  /* <dr2> */  input arx_17_h,
  /* <dl2> */  input arx_18_a_h,
  /* <cp1> */  input arx_19_a_h,
  /* <cm1> */  input arx_20_h,
  /* <ck2> */  input arx_21_h,
  /* <cf1> */  input arx_22_h,
  /* <ck1> */  input arx_23_h,
  /* <cf2> */  input arx_24_a_h,
  /* <cd1> */  input arx_25_a_h,
  /* <dd2> */  input arx_26_h,
  /* <de2> */  input arx_27_h,
  /* <fd2> */  input arx_28_h,
  /* <fa1> */  input arx_29_h,
  /* <fl1> */  input arx_30_a_h,
  /* <fe1> */  input arx_31_a_h,
  /* <ed2> */  input arx_32_h,
  /* <dp1> */  input arx_33_h,
  /* <dj2> */  input arx_34_h,
  /* <dk2> */  input arx_35_h,
  /* <et2> */  input con_ar_36_h,
  /* <fn1> */  input con_arx_36_h,
  /* <de1> */  input cram_shNgarmm_sel_1_a_h,
  /* <da1> */  input cram_shNgarmm_sel_2_a_h,
  /* <dm1> */  input scd2_sc_04_h,
  /* <dk1> */  input scd2_sc_05_h,
  /* <dj1> */  input scd2_sc_06_h,
  /* <df1> */  input scd2_sc_07_h,
  /* <cp2> */  input scd2_sc_08_h,
  /* <cs2> */  input scd2_sc_09_h,
  /* <ch2> */  input scd2_sc_36_to_63_h,
  /* <dd1> */  input scd2_sc_DtgeDt_36_h,
  /* <bl1> */ output sh_00_h,
  /* <bk1> */ output sh_01_h,
  /* <bj1> */ output sh_02_h,
  /* <bf1> */ output sh_03_h,
  /* <af2> */ output sh_04_h,
  /* <ae2> */ output sh_05_h,
  /* <af1> */ output sh_06_h,
  /* <ae1> */ output sh_07_h,
  /* <am2> */ output sh_08_h,
  /* <am1> */ output sh_09_h,
  /* <ba1> */ output sh_10_h,
  /* <av2> */ output sh_11_h,
  /* <bk2> */ output sh_12_h,
  /* <bf2> */ output sh_13_h,
  /* <bd2> */ output sh_14_h,
  /* <as2> */ output sh_15_h,
  /* <ap2> */ output sh_16_h,
  /* <al1> */ output sh_17_h,
  /* <aj2> */ output sh_18_h,
  /* <ad2> */ output sh_19_h,
  /* <aj1> */ output sh_20_h,
  /* <ad1> */ output sh_21_h,
  /* <ak2> */ output sh_22_h,
  /* <aa1> */ output sh_23_h,
  /* <ar2> */ output sh_24_h,
  /* <ak1> */ output sh_25_h,
  /* <au2> */ output sh_26_h,
  /* <ar1> */ output sh_27_h,
  /* <bp2> */ output sh_28_h,
  /* <bl2> */ output sh_29_h,
  /* <bm2> */ output sh_30_h,
  /* <bj2> */ output sh_31_h,
  /* <be2> */ output sh_32_h,
  /* <as1> */ output sh_33_h,
  /* <ap1> */ output sh_34_h,
  /* <al2> */ output sh_35_h,
  /* <cs1> */ output sh_ar_par_odd_a_h,
  /* <dc1> */ output shm1_ar_extended_h,
  /* <cu2> */ output shm1_ar_par_odd_a_l,
  /* <ed1> */ output shm1_ar_par_odd_b_h,
  /* <ea1> */ output shm1_ar_par_odd_b_l,
  /* <cv2> */ output shm1_ar_par_odd_h,
  /* <fe2> */ output shm1_arx_par_odd_h,
  /* <dr1> */ output shm1_indexed_h,
  /* <ds1> */ output shm1_xr_01_h,
  /* <dh2> */ output shm1_xr_02_h,
  /* <ec1> */ output shm1_xr_04_h,
  /* <dt2> */ output shm1_xr_10_h,
  /* <bp1> */ output shm4_sh_00_a_h,
  /* <bm1> */ output shm4_sh_01_a_h,
  /* <be1> */ output shm4_sh_02_a_h,
  /* <bd1> */ output shm4_sh_03_a_h
);

`include "shm46.svh"

endmodule	// shm46
