module mbc22(
  /* <ev2> */ output a_change_coming_in_l,
  /* <er1> */ output ackn_pulse_l,
  /* <es1> */  input apr2_wr_bad_adr_par_l,
  /* <aj2> */ output cache_adr_27_h,
  /* <ak1> */ output cache_adr_28_h,
  /* <ak2> */ output cache_adr_29_h,
  /* <am2> */ output cache_adr_30_h,
  /* <aa1> */ output cache_adr_31_h,
  /* <ac1> */ output cache_adr_32_h,
  /* <ad2> */ output cache_adr_33_h,
  /* <cf1> */ output cache_adr_34_h,
  /* <da1> */ output cache_adr_35_h,
  /* <cm2> */ output cache_adr_35_l,
  /* <cl2> */ output cache_wr_00_a_l,
  /* <ck1> */ output cache_wr_09_a_l,
  /* <ch2> */ output cache_wr_18_a_l,
  /* <cj2> */ output cache_wr_27_a_l,
  /* <cs2> */ output cam_sel_1_h,
  /* <bj2> */ output cam_sel_2_h,
  /* <df2> */  input ccl_start_mem_l,
  /* <cr2> */  input clk1_mbc_h,
  /* <ee1> */ output core_busy_a_h,
  /* <ds1> */  input core_busy_h,
  /* <ef1> */ output core_rd_in_prog_h,
  /* <dl2> */  input csh2_e_core_rd_rq_b_l,
  /* <et2> */  input csh2_one_word_rd_h,
  /* <el1> */  input csh2_rd_pause_2nd_half_l,
  /* <am1> */  input csh3_adr_pma_en_h,
  /* <df1> */  input csh3_any_val_hold_a_h,
  /* <bf1> */  input csh3_match_hold_1_in_h,
  /* <be2> */  input csh3_match_hold_2_in_h,
  /* <dl1> */  input csh4_clear_wr_t0_l,
  /* <es2> */  input csh4_data_clr_done_l,
  /* <dm2> */  input csh4_ebox_t3_l,
  /* <fn1> */  input csh4_ebox_wr_t4_in_h,
  /* <cr1> */  input csh5_chan_rd_t5_l,
  /* <dr1> */  input csh5_chan_t3_l,
  /* <fr2> */  input csh5_chan_wr_t5_in_h,
  /* <de1> */  input csh5_page_refill_t9_l,
  /* <fl2> */  input csh6_cache_wr_in_h,
  /* <ep1> */  input csh6_chan_wr_cache_l,
  /* <fm2> */  input csh6_wr_from_mem_nxt_h,
  /* <br1> */ output csh_0_wr_en_l,
  /* <bd1> */ output csh_1_wr_en_l,
  /* <dc1> */ output csh_2_wr_en_l,
  /* <cf2> */ output csh_3_wr_en_l,
  /* <fl1> */ output csh_adr_wr_pulse_l,
  /* <cp2> */ output csh_sel_lru_h,
  /* <dm1> */ output csh_sel_lru_l,
  /* <cd2> */ output csh_val_sel_all_h,
  /* <cn1> */ output csh_val_wr_data_h,
  /* <fp1> */ output csh_val_wr_pulse_l,
  /* <dj2> */ output csh_wr_sel_all_h,
  /* <ek2> */ output csh_wr_wr_data_h,
  /* <fp2> */ output csh_wr_wr_pulse_l,
  /* <br2> */ output data_valid_a_out_h,
  /* <dh2> */ output data_valid_b_out_h,
  /* <bc1> */  input diag_04_b_h,
  /* <ba1> */  input diag_05_b_h,
  /* <au2> */  input diag_06_b_h,
  /* <at2> */  input diag_read_func_16x_l,
  /* <eu2> */  input e_cache_wr_cyc_l,
  /* <cj1> */ output ebus_d27_e_h,
  /* <cl1> */ output ebus_d28_e_h,
  /* <ct2> */ output ebus_d29_e_h,
  /* <dd1> */ output ebus_d30_e_h,
  /* <dd2> */ output ebus_d31_e_h,
  /* <dj1> */ output ebus_d32_e_h,
  /* <dk1> */ output ebus_d33_e_h,
  /* <cu2> */  input force_valid_match_0_h,
  /* <bm1> */  input force_valid_match_1_h,
  /* <ca1> */  input force_valid_match_2_h,
  /* <cm1> */  input force_valid_match_3_h,
  /* <ae2> */  input load_ebus_reg_l,
  /* <bs1> */  input mb_sel_1_h,
  /* <ce1> */  input mb_sel_2_h,
  /* <ee2> */ output mbc1_write_ok_h,
  /* <cv2> */ output mbc2_csh_data_clr_t1_l,
  /* <bm2> */ output mbc2_csh_data_clr_t2_l,
  /* <cc1> */ output mbc2_csh_data_clr_t3_l,
  /* <bp2> */ output mbc2_data_clr_done_in_l,
  /* <ef2> */ output mbc3_a_change_coming_a_l,
  /* <dk2> */ output mbc3_a_phase_coming_l,
  /* <em2> */ output mbc3_csh_wr_wr_data_l,
  /* <bj1> */ output mbc3_inh_1st_mb_req_h,
  /* <ej2> */ output mbc4_core_adr_34_h,
  /* <bf2> */ output mbc4_core_adr_35_h,
  /* <bt2> */ output mbc4_core_data_val_Ng1_l,
  /* <ep2> */ output mbc4_core_data_val_Ng2_l,
  /* <ff2> */ output mbc4_core_data_valid_h,
  /* <fr1> */ output mbc4_core_data_valid_l,
  /* <dv2> */ output mbc4_mem_start_l,
  /* <fm1> */  input mbx1_cca_inval_t4_a_h,
  /* <aj1> */  input mbx1_refill_adr_en_h,
  /* <dp2> */  input mbx2_chan_wr_cyc_l,
  /* <cd1> */  input mbx3_refill_hold_h,
  /* <em1> */  input mbx4_cache_to_mb_t2_l,
  /* <dn1> */  input mbx4_cache_to_mb_t4_a_l,
  /* <fs1> */  input mbx4_writeback_t2_h,
  /* <fe1> */  input mbx5_mem_rd_rq_in_h,
  /* <fc1> */  input mbx5_mem_to_c_en_l,
  /* <fv2> */  input mbx5_rq_0_in_h,
  /* <fn2> */  input mbx5_rq_0_in_h,
  /* <fu2> */  input mbx5_rq_1_in_h,
  /* <ft2> */  input mbx5_rq_2_in_h,
  /* <fs2> */  input mbx5_rq_3_in_h,
  /* <av2> */ output mbx_csh_adr_27_h,
  /* <ap2> */ output mbx_csh_adr_28_h,
  /* <ar2> */ output mbx_csh_adr_29_h,
  /* <an1> */ output mbx_csh_adr_30_h,
  /* <al1> */ output mbx_csh_adr_31_h,
  /* <af2> */ output mbx_csh_adr_32_h,
  /* <ad1> */ output mbx_csh_adr_33_h,
  /* <ed2> */  input mem_ackn_a_h,
  /* <ed1> */  input mem_ackn_b_h,
  /* <bh2> */ output mem_adr_par_h,
  /* <ea1> */  input mem_data_valid_a_l,
  /* <ec1> */  input mem_data_valid_b_l,
  /* <cs1> */ output mem_rd_rq_b_h,
  /* <ej1> */ output mem_rd_rq_h,
  /* <bk2> */ output mem_rq_0_h,
  /* <bu2> */ output mem_rq_1_h,
  /* <ck2> */ output mem_rq_2_h,
  /* <du2> */ output mem_rq_3_h,
  /* <dr2> */ output mem_start_a_h,
  /* <dp1> */ output mem_start_b_h,
  /* <bs2> */ output mem_to_c_en_l,
  /* <eh2> */ output mem_wr_rq_h,
  /* <bl2> */ output mem_wr_rq_l,
  /* <ce2> */  input mr_reset_06_h,
  /* <er2> */  input nxm_ackn_h,
  /* <fe2> */  input nxm_data_val_l,
  /* <en1> */ output phase_change_coming_l,
  /* <bd2> */  input pma3_pa_27_h,
  /* <ar1> */  input pma3_pa_28_h,
  /* <as2> */  input pma3_pa_29_h,
  /* <af1> */  input pma3_pa_30_h,
  /* <al2> */  input pma3_pa_31_h,
  /* <cp1> */  input pma4_34_b_h,
  /* <de2> */  input pma4_35_b_h,
  /* <fk2> */  input pma4_adr_par_h,
  /* <ah2> */  input pma4_pa_32_h,
  /* <ae1> */  input pma4_pa_33_h,
  /* <ds2> */  input pma5_csh_writeback_cyc_l,
  /* <bp1> */ output rq_hold_ff_h,
  /* <fj2> */  input sbus_adr_34_h,
  /* <fj1> */  input sbus_adr_35_h,
  /* <dt2> */ output sbus_adr_hold_h
);

`include "mbc22.svh"

endmodule	// mbc22
