module just_a_wire(input bit b, output bit q);
  always_comb q = b;
endmodule // just_a_wire
