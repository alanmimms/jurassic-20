module pag;
`include "pag.svh"
endmodule	// pag
