module clk;
`include "clk.svh"
endmodule	// clk
