module mtr33(
  /* <es2> */ input  ch_t1_h,
  /* <ep2> */ input  chc1_cbus_ready_e_l,
  /* <cr2> */ input  clk1_mtr_h,
  /* <aj2> */ input  clk3_ebox_sync_c_l,
  /* <du2> */ input  clk_mb_xfer_l,
  /* <da1> */ input  con_mbox_wait_l,
  /* <cj2> */ input  con_pi_cycle_b_h,
  /* <dk2> */ input  con_ucode_state_01_h,
  /* <dc1> */ input  con_ucode_state_03_h,
  /* <ae2> */ input  cram_Nr_06_a_h,
  /* <ad2> */ input  cram_Nr_07_a_h,
  /* <ah2> */ input  cram_Nr_08_a_h,
  /* <em2> */ input  crc_sel_1d_l,
  /* <ej2> */ input  crc_sel_2d_l,
  /* <eh2> */ input  crc_sel_4d_l,
  /* <fk2> */ input  csh7_cca_writeback_l,
  /* <fm2> */ output csh7_cca_writeback_l,
  /* <fp2> */ input  csh7_e_writeback_l,
  /* <ft2> */ input  csh7_e_writeback_l,
  /* <fv2> */ input  csh7_fill_cache_rd_l,
  /* <fs2> */ input  csh7_fill_cache_rd_l,
  /* <af2> */ input  ctl1_spec_mtr_ctl_l,
  /* <ct2> */ input  ctl3_diag_rd_func_11x_l,
  /* <de2> */ input  diag_04_b_h,
  /* <df2> */ input  diag_05_b_h,
  /* <dd2> */ input  diag_06_b_h,
  /* <bl2> */ input  ebus_d18_e_h,
  /* <bk2> */ input  ebus_d19_e_h,
  /* <bm2> */ output ebus_d20_e_h,
  /* <be2> */ output ebus_d21_e_h,
  /* <bf2> */ output ebus_d22_e_h,
  /* <bd2> */ output ebus_d23_e_h,
  /* <dm1> */ output ebus_d24_e_h,
  /* <dn1> */ output ebus_d25_e_h,
  /* <dl1> */ output ebus_d26_e_h,
  /* <dj1> */ output ebus_d27_e_h,
  /* <dj2> */ output ebus_d28_e_h,
  /* <dk1> */ output ebus_d29_e_h,
  /* <fa1> */ output ebus_d30_e_h,
  /* <fk1> */ output ebus_d31_e_h,
  /* <fc1> */ output ebus_d32_e_h,
  /* <fh2> */ output ebus_d33_e_h,
  /* <fe2> */ output ebus_d34_e_h,
  /* <fj1> */ output ebus_d35_e_h,
  /* <dh2> */ input  mr_reset_02_h,
  /* <dl2> */ input  mtr1_cache_cry_10_in_l,
  /* <dm2> */ output mtr1_cache_cry_10_l,
  /* <dr1> */ input  mtr1_ebox_cry_10_in_l,
  /* <dp2> */ output mtr1_ebox_cry_10_l,
  /* <fr1> */ input  mtr1_interval_cry_14_in_l,
  /* <fs1> */ output mtr1_interval_cry_14_l,
  /* <cd2> */ input  mtr1_perf_cry_10_in_l,
  /* <ce2> */ output mtr1_perf_cry_10_l,
  /* <dt2> */ input  mtr1_time_cry_10_in_l,
  /* <dv2> */ output mtr1_time_cry_10_l,
  /* <fr2> */ output mtr4_e_writeback_l,
  /* <fu2> */ output mtr4_fill_cache_rd_l,
  /* <ed2> */ output mtr_1_mhz_a_l,
  /* <fl2> */ input  mtr_cca_writeback_l,
  /* <as2> */ output mtr_cono_mtrCm_l,
  /* <at2> */ output mtr_interrupt_req_h,
  /* <ak2> */ output mtr_vector_interrupt_l,
  /* <ch2> */ input  pi2_hold_1_h,
  /* <cp2> */ input  pi2_hold_2_h,
  /* <ck2> */ input  pi2_hold_4_h,
  /* <cf2> */ input  pi2_pi1_a_h,
  /* <cl2> */ input  pi2_pi2_a_h,
  /* <cm2> */ input  pi2_pi4_a_h,
  /* <fd2> */ input  pi3_mtr_pia_01_h,
  /* <ff2> */ input  pi3_mtr_pia_02_h,
  /* <fj2> */ input  pi3_mtr_pia_04_h,
  /* <ca1> */ input  probe_h,
  /* <cu2> */ input  scd_user_a_l,
  /* <cc1> */ input  vma1_ac_ref_a_l
);

`include "mtr33nets.svh"

endmodule	// mtr33
