module top(input clk60);

   

endmodule // top
