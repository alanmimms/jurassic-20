module crc10(
  /* <dh2> */  input ccl_act_flag_req_l,
  /* <cj1> */  input ccl_ccwf_clr_h,
  /* <bp2> */  input ccl_error_h,
  /* <ef2> */  input ccl_last_xfer_err_in_h,
  /* <br2> */  input ccl_load_ac_h,
  /* <bm2> */  input ccl_load_ac_l,
  /* <ae2> */  input ccl_mb_cyc_t2_l,
  /* <dj2> */  input ccl_mb_req_t2_l,
  /* <dd2> */  input ccl_mem_store_req_l,
  /* <ej2> */  input ccl_op_load_h,
  /* <ef1> */  input ccl_op_load_l,
  /* <at2> */  input ccl_ram_req_l,
  /* <ad2> */  input ccl_req_ctr_en_l,
  /* <ct2> */  input ccl_wcEq0_in_h,
  /* <df2> */  input ccl_wcEq0_in_l,
  /* <bl2> */  input ccw_act_ctr_0_en_l,
  /* <be2> */  input ccw_act_ctr_1_en_l,
  /* <bf2> */  input ccw_act_ctr_2_en_l,
  /* <ep2> */  input ccw_buf_00_in_l,
  /* <en1> */  input ccw_buf_01_in_l,
  /* <eh2> */  input ccw_buf_02_in_l,
  /* <ch2> */  input ccw_ccwf_waiting_h,
  /* <av2> */  input ch_cbus_req_h,
  /* <ds2> */  input ch_cbus_req_l,
  /* <au2> */  input ch_contr_req_h,
  /* <cf2> */  input ch_contr_req_l,
  /* <ep1> */  input ch_done_intr_l,
  /* <bt2> */  input ch_mr_reset_b_h,
  /* <ff2> */  input ch_req_d_l,
  /* <cv2> */  input ch_reset_intr_h,
  /* <el1> */  input ch_reset_intr_l,
  /* <cu2> */  input ch_start_intr_h,
  /* <ck2> */  input ch_start_intr_l,
  /* <cl2> */  input ch_start_l,
  /* <du2> */  input ch_store_h,
  /* <cr2> */  input clk_crc_h,
  /* <bh2> */ output crc_act_ctr_0_h,
  /* <bj2> */ output crc_act_ctr_1_h,
  /* <bd2> */ output crc_act_ctr_2_h,
  /* <bk2> */ output crc_act_ctr_2r_l,
  /* <de2> */ output crc_act_flag_ena_l,
  /* <fr1> */ output crc_cbus_contr_cyc_l,
  /* <ee1> */ output crc_cbus_out_hold_h,
  /* <cj2> */ output crc_ccwf_en_l,
  /* <ev2> */ output crc_err_in_h,
  /* <ed2> */ output crc_last_word_in_h,
  /* <em2> */ output crc_long_wc_err_h,
  /* <ek1> */ output crc_mb_cyc_h,
  /* <fn1> */ output crc_mb_cyc_l,
  /* <ed1> */ output crc_mem_store_ena_l,
  /* <el2> */ output crc_ovn_err_in_h,
  /* <as2> */  input crc_ram_adr_1r_h,
  /* <ar2> */  input crc_ram_adr_2r_h,
  /* <am2> */  input crc_ram_adr_4r_h,
  /* <cs2> */ output crc_ram_cyc_l,
  /* <dr1> */ output crc_ready_in_h,
  /* <dt2> */ output crc_req_d_h,
  /* <fv2> */ output crc_req_e_l,
  /* <ek2> */ output crc_reset_l,
  /* <em1> */ output crc_reverse_in_h,
  /* <dr2> */ output crc_rh20_err_in_h,
  /* <eu2> */ output crc_short_wc_err_h,
  /* <ap2> */  input crc_wr_ram_l
);

`include "crc10nets.svh"

endmodule	// crc10
