module con35(
  /* <fp1> */  input apr_fm_36_h,
  /* <cr2> */  input clk_con_h,
  /* <ba1> */  input clk_ebox_sync_a_l,
  /* <fk1> */  input clk_mb_xfer_h,
  /* <ap1> */  input clk_page_error_h,
  /* <fn1> */  input clk_sbr_call_h,
  /* <ck2> */ output con1_condSl024_l,
  /* <dm1> */ output con2_long_en_l,
  /* <be2> */ output con3_Nr_func_010_h,
  /* <bd1> */ output con3_Nr_func_011_h,
  /* <ek1> */ output con3_Nr_func_04x_l,
  /* <ek2> */ output con3_Nr_func_05x_l,
  /* <fd2> */ output con4_spec_08_h,
  /* <ak2> */ output con_ar_36_h,
  /* <ev2> */ output con_ar_36_l,
  /* <ef1> */ output con_ar_from_ebus_h,
  /* <el2> */ output con_ar_loaded_l,
  /* <aj2> */ output con_arx_36_h,
  /* <ej1> */ output con_arx_loaded_l,
  /* <ar1> */ output con_cache_load_en_h,
  /* <ae1> */ output con_cache_look_en_l,
  /* <bk1> */ output con_clr_private_instr_h,
  /* <cj1> */ output con_condSl026_l,
  /* <cj2> */ output con_condSl027_l,
  /* <ce1> */ output con_condSlad_flags_h,
  /* <ee1> */ output con_condSldiag_func_l,
  /* <du2> */ output con_condSlebus_ctl_l,
  /* <cf2> */ output con_condSlfe_shrt_h,
  /* <cn1> */ output con_condSlload_vma_held_h,
  /* <cp1> */ output con_condSlmbox_ctl_l,
  /* <cf1> */ output con_condSlpcfGETSNr_h,
  /* <cd1> */ output con_condSlsel_vma_h,
  /* <cp2> */ output con_condSlsel_vma_l,
  /* <ct2> */ output con_condSlvmaGETSNr_h,
  /* <bm2> */ output con_cond_adr_10_h,
  /* <cm2> */ output con_cond_en_00to07_l,
  /* <cm1> */ output con_cond_en_30to37_l,
  /* <dc1> */ output con_cond_instr_abort_h,
  /* <fv2> */ output con_cono_200000_h,
  /* <dd1> */ output con_cono_apr_l,
  /* <aj1> */ output con_cono_pi_l,
  /* <as2> */ output con_datao_apr_l,
  /* <al2> */ output con_delay_req_h,
  /* <en1> */ output con_ebox_halted_h,
  /* <bt2> */ output con_ebus_rel_h,
  /* <fe1> */ output con_fm_write_00to17_l,
  /* <ed1> */ output con_fm_write_18to35_l,
  /* <ff1> */ output con_fm_write_par_l,
  /* <fl1> */ output con_fm_xfer_h,
  /* <fj1> */ output con_fm_xfer_l,
  /* <aa1> */ output con_ki10_paging_mode_h,
  /* <bl2> */ output con_ki10_paging_mode_l,
  /* <ej2> */ output con_load_ac_blocks_l,
  /* <br2> */ output con_load_access_cond_h,
  /* <bp2> */ output con_load_dram_h,
  /* <eu2> */ output con_load_dram_l,
  /* <bs2> */ output con_load_ir_l,
  /* <eh2> */ output con_load_prev_context_l,
  /* <et2> */ output con_load_spec_instr_l,
  /* <fh2> */ output con_mbox_wait_l,
  /* <bj1> */ output con_nicond_07_h,
  /* <bh2> */ output con_nicond_08_h,
  /* <bf1> */ output con_nicond_09_h,
  /* <bj2> */ output con_nicond_trap_en_h,
  /* <fa1> */ output con_pcPl1_inh_h,
  /* <bk2> */ output con_pcPl1_inh_l,
  /* <es1> */ output con_pi_cycle_a_h,
  /* <es2> */ output con_pi_cycle_a_l,
  /* <ep2> */ output con_pi_cycle_b_h,
  /* <er2> */ output con_pi_cycle_b_l,
  /* <er1> */ output con_pi_disable_l,
  /* <fk2> */ output con_pi_dismiss_l,
  /* <bs1> */ output con_run_h,
  /* <de1> */ output con_sel_clr_h,
  /* <dh2> */ output con_sel_dis_h,
  /* <df2> */ output con_sel_en_l,
  /* <dd2> */ output con_sel_set_l,
  /* <fe2> */ output con_set_pih_l,
  /* <cl2> */ output con_skip_en_40to47_l,
  /* <ck1> */ output con_skip_en_50to57_l,
  /* <be1> */ output con_sr_00_h,
  /* <cr1> */ output con_sr_01_h,
  /* <cs1> */ output con_sr_02_h,
  /* <cs2> */ output con_sr_03_h,
  /* <ac1> */ output con_trap_en_a_h,
  /* <da1> */ output con_trap_en_h,
  /* <ef2> */ output con_ucode_state_01_h,
  /* <ee2> */ output con_ucode_state_03_h,
  /* <ed2> */ output con_ucode_state_07_h,
  /* <ar2> */ output con_vma_sel_1_l,
  /* <an1> */ output con_vma_sel_2_l,
  /* <am2> */ output con_wr_even_par_adr_h,
  /* <af2> */ output con_wr_even_par_dir_l,
  /* <ec1> */  input cram_Nr_00_e_h,
  /* <ea1> */  input cram_Nr_01_e_h,
  /* <el1> */  input cram_Nr_02_e_h,
  /* <dt2> */  input cram_Nr_03_e_h,
  /* <dn1> */  input cram_Nr_04_e_h,
  /* <em1> */  input cram_Nr_05_e_h,
  /* <dk1> */  input cram_Nr_06_e_h,
  /* <bc1> */  input cram_Nr_07_e_h,
  /* <dp1> */  input cram_Nr_08_e_h,
  /* <ah2> */  input cram_cond_00_h,
  /* <af1> */  input cram_cond_01_h,
  /* <ak1> */  input cram_cond_02_h,
  /* <ad2> */  input cram_cond_03_h,
  /* <ad1> */  input cram_cond_04_h,
  /* <ae2> */  input cram_cond_05_h,
  /* <fl2> */  input cram_mem_02_a_l,
  /* <fr1> */  input csh_par_bit_a_h,
  /* <fp2> */  input csh_par_bit_b_h,
  /* <em2> */  input ctl_console_control_h,
  /* <dj2> */  input ctl_dispSlnicond_h,
  /* <fm1> */  input ctl_ebus_xfer_l,
  /* <fd1> */  input ctl_specSlflag_ctl_l,
  /* <fc1> */  input ctl_specSlsave_flags_l,
  /* <at2> */  input diag_06_a_h,
  /* <ds2> */  input diag_control_func_01x_l,
  /* <ca1> */ output ebus_d18_e_h,
  /* <cd2> */ output ebus_d19_e_h,
  /* <ce2> */ output ebus_d20_e_h,
  /* <cc1> */ output ebus_d21_e_h,
  /* <cu2> */ output ebus_d22_e_h,
  /* <cv2> */ output ebus_d23_e_h,
  /* <dv2> */ output ebus_d24_e_h,
  /* <dr1> */  input ebus_ds04_e_h,
  /* <dp2> */  input ebus_ds05_e_h,
  /* <dr2> */  input ebus_ds06_e_h,
  /* <fu2> */  input ebus_parity_active_e_h,
  /* <fm2> */  input ebus_parity_e_h,
  /* <ds1> */  input ir_IO_legal_h,
  /* <ap2> */  input mbz1_rdNgpseNgwr_ref_l,
  /* <ft2> */  input mcl_load_ar_h,
  /* <al1> */  input mcl_load_vma_h,
  /* <ep1> */  input mcl_mbox_cyc_req_h,
  /* <ff2> */  input mcl_skip_satisfied_h,
  /* <fr2> */  input mcl_store_ar_l,
  /* <fs2> */  input mcl_vma_fetch_l,
  /* <cl1> */  input mcl_vma_section_0_h,
  /* <df1> */  input mr_reset_04_h,
  /* <dk2> */  input mtr_interrupt_req_h,
  /* <bu2> */  input pi2_ext_tran_rec_h,
  /* <dj1> */  input pi2_ready_h,
  /* <bv2> */  input pi5_ebus_cp_grant_h,
  /* <as1> */  input scd_public_a_l,
  /* <dl2> */  input scd_user_a_l,
  /* <dl1> */  input scd_user_iot_a_l,
  /* <de2> */  input vma_ac_ref_l
);

`include "con35nets.svh"

endmodule	// con35
