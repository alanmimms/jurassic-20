module scd;
`include "scd.svh"
endmodule	// scd
