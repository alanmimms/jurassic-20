module cra;
`include "cra.svh"
endmodule	// cra
