module csh23(
  /* <bc1> */ input  a_change_coming_in_l,
  /* <da1> */ input  apr6_ebox_cca_l,
  /* <ba1> */ input  apr6_ebox_era_l,
  /* <ds1> */ input  apr6_ebox_load_reg_l,
  /* <aj1> */ input  apr6_ebox_read_reg_h,
  /* <av2> */ input  apr6_ebox_read_reg_l,
  /* <ak1> */ input  apr6_ebox_sbus_diag_h,
  /* <dk1> */ input  apr_ebox_sbus_diag_l,
  /* <fr1> */ input  apr_en_refill_ram_wr_h,
  /* <ef2> */ input  cache_to_mb_t4_l,
  /* <fe1> */ input  ccl_chan_req_h,
  /* <fl1> */ input  ccl_chan_req_l,
  /* <af1> */ input  ccl_chan_to_mem_h,
  /* <dt2> */ input  ccl_chan_to_mem_l,
  /* <ce1> */ input  chan_read_h,
  /* <cr2> */ input  clk1_csh_h,
  /* <ej2> */ input  clk3_ebox_sync_d_l,
  /* <fa1> */ input  clk4_ebox_cyc_abort_h,
  /* <fh2> */ input  clk4_ebox_req_h,
  /* <ee1> */ input  clk4_ebox_req_l,
  /* <at2> */ input  con_ki10_paging_mode_h,
  /* <ec1> */ input  core_busy_h,
  /* <fv2> */ input  core_busy_l,
  /* <ap2> */ output csh1_cca_cyc_l,
  /* <eu2> */ output csh1_cca_req_grant_h,
  /* <ev2> */ output csh1_chan_req_grant_h,
  /* <ca1> */ output csh1_ebox_cca_grant_h,
  /* <aa1> */ output csh1_ebox_era_grant_h,
  /* <es1> */ output csh1_ebox_req_grant_a_l,
  /* <ek2> */ output csh1_ebox_req_grant_h,
  /* <bp2> */ output csh1_mb_cyc_l,
  /* <et2> */ output csh1_mb_req_grant_l,
  /* <bk2> */ output csh1_pgrf_cyc_a_h,
  /* <bj2> */ output csh1_pgrf_cyc_a_l,
  /* <fm1> */ output csh1_ready_to_go_h,
  /* <cc1> */ output csh1_ready_to_go_l,
  /* <em2> */ output csh2_e_cache_wr_cyc_h,
  /* <ea1> */ output csh2_e_core_rd_rq_b_l,
  /* <fs2> */ output csh2_e_core_rd_rq_l,
  /* <as1> */ output csh2_ebox_retry_req_l,
  /* <bd1> */ output csh2_mbox_resp_in_h,
  /* <bk1> */ output csh2_one_word_rd_h,
  /* <be2> */ output csh2_one_word_rd_l,
  /* <dp2> */ output csh2_rd_pause_2nd_half_l,
  /* <ep2> */ output csh3_adr_pma_en_h,
  /* <fj1> */ output csh3_adr_ready_l,
  /* <fr2> */ output csh3_any_val_hold_a_h,
  /* <ff1> */ output csh3_any_val_hold_in_h,
  /* <ep1> */ output csh3_gate_vma_27to33_h,
  /* <br2> */ output csh3_match_hold_1_in_h,
  /* <bu2> */ output csh3_match_hold_2_in_h,
  /* <fm2> */ output csh3_mb_wr_rq_clr_nxt_l,
  /* <ck1> */ output csh4_clear_wr_t0_l,
  /* <er2> */ output csh4_data_clr_done_l,
  /* <fd1> */ output csh4_ebox_t0_in_h,
  /* <au2> */ output csh4_ebox_t3_l,
  /* <dh2> */ output csh4_ebox_wr_t4_in_h,
  /* <dj1> */ output csh4_one_word_wr_t0_l,
  /* <fs1> */ output csh4_writeback_t1_a_l,
  /* <ee2> */ output csh5_chan_rd_t5_l,
  /* <ad1> */ output csh5_chan_t3_l,
  /* <ds2> */ output csh5_chan_t4_l,
  /* <dr2> */ output csh5_chan_wr_t5_in_h,
  /* <bt2> */ output csh5_page_refill_t12_l,
  /* <dj2> */ output csh5_page_refill_t4_l,
  /* <ar2> */ output csh5_page_refill_t8_l,
  /* <cj1> */ output csh5_page_refill_t9_l,
  /* <em1> */ output csh5_t2_l,
  /* <am2> */ output csh6_cache_wr_in_h,
  /* <dm2> */ output csh6_cca_cyc_done_l,
  /* <ap1> */ output csh6_cca_inval_t4_l,
  /* <ad2> */ output csh6_chan_wr_cache_l,
  /* <cn1> */ output csh6_ebox_load_reg_h,
  /* <cd2> */ output csh6_mbox_pt_dir_wr_l,
  /* <cf2> */ output csh6_page_fail_hold_h,
  /* <df2> */ output csh6_page_fail_hold_l,
  /* <bp1> */ output csh6_page_refill_error_h,
  /* <bm1> */ output csh6_page_refill_error_l,
  /* <fp1> */ output csh6_wr_from_mem_nxt_h,
  /* <el1> */ output csh7_cca_writeback_l,
  /* <fk1> */ output csh7_e_writeback_l,
  /* <ft2> */ output csh7_fill_cache_rd_l,
  /* <ck2> */ input  csh_0_any_wr_l,
  /* <bj1> */ input  csh_0_valid_match_h,
  /* <cu2> */ input  csh_0_valid_match_l,
  /* <de2> */ input  csh_0_wd_val_h,
  /* <cm2> */ input  csh_1_any_wr_l,
  /* <bs2> */ input  csh_1_valid_match_h,
  /* <cv2> */ input  csh_1_valid_match_l,
  /* <df1> */ input  csh_1_wd_val_h,
  /* <cl2> */ input  csh_2_any_wr_l,
  /* <bv2> */ input  csh_2_valid_match_h,
  /* <ct2> */ input  csh_2_valid_match_l,
  /* <dc1> */ input  csh_2_wd_val_h,
  /* <cp1> */ input  csh_3_any_wr_l,
  /* <bs1> */ input  csh_3_valid_match_h,
  /* <cs2> */ input  csh_3_valid_match_l,
  /* <dd2> */ input  csh_3_wd_val_h,
  /* <ak2> */ output csh_chan_cyc_l,
  /* <du2> */ output csh_ebox_cyc_a_l,
  /* <cr1> */ input  csh_lru_1_h,
  /* <cj2> */ input  csh_lru_2_h,
  /* <fl2> */ output csh_refill_ram_wr_l,
  /* <es2> */ output csh_use_hold_h,
  /* <ar1> */ output csh_use_wr_en_h,
  /* <dl2> */ input  ctl3_diag_ld_ebus_reg_l,
  /* <dp1> */ input  diag_04_b_h,
  /* <dr1> */ input  diag_05_b_h,
  /* <dm1> */ input  diag_06_b_h,
  /* <ef1> */ input  diag_read_func_17x_l,
  /* <bh2> */ output e_cache_wr_cyc_l,
  /* <al1> */ output ebus_d22_e_h,
  /* <am1> */ output ebus_d23_e_h,
  /* <cd1> */ output ebus_d24_e_h,
  /* <cm1> */ output ebus_d25_e_h,
  /* <fd2> */ output ebus_d26_e_h,
  /* <el2> */ output ebus_d27_e_h,
  /* <er1> */ output ebus_d28_e_h,
  /* <dk2> */ output ebus_d29_e_h,
  /* <br1> */ output load_ebus_reg_l,
  /* <cf1> */ output mb_test_par_a_in_l,
  /* <dd1> */ input  mbc1_write_ok_h,
  /* <af2> */ input  mbc2_csh_data_clr_t1_l,
  /* <bf1> */ input  mbc2_csh_data_clr_t2_l,
  /* <ek1> */ input  mbc2_csh_data_clr_t3_l,
  /* <eh2> */ input  mbc2_data_clr_done_in_l,
  /* <bl1> */ input  mbc4_core_data_val_Ng1_l,
  /* <ae1> */ input  mbc4_core_data_valid_h,
  /* <be1> */ input  mbc4_core_data_valid_l,
  /* <ah2> */ input  mbx1_cache_bit_h,
  /* <ce2> */ input  mbx1_cache_bit_l,
  /* <bf2> */ input  mbx1_cca_all_pages_cyc_l,
  /* <al2> */ input  mbx1_csh_cca_inval_csh_h,
  /* <aj2> */ input  mbx1_csh_cca_val_core_h,
  /* <ac1> */ input  mbx1_csh_cca_val_core_l,
  /* <fc1> */ input  mbx1_refill_adr_en_nxt_h,
  /* <fu2> */ input  mbx2_mb_sel_hold_ff_h,
  /* <cp2> */ input  mbx2_mb_sel_hold_l,
  /* <bd2> */ input  mbx3_sbus_diag_3_l,
  /* <fk2> */ input  mbx4_cache_to_mb_done_l,
  /* <cs1> */ input  mbx5_mb_req_in_h,
  /* <ej1> */ input  mcl2_vma_pause_h,
  /* <fj2> */ input  mcl2_vma_read_l,
  /* <dv2> */ input  mcl2_vma_write_l,
  /* <cl1> */ input  mcl6_ebox_map_l,
  /* <bl2> */ input  mem_busy_h,
  /* <ae2> */ input  mr_reset_05_h,
  /* <as2> */ input  pag4_page_fail_l,
  /* <ed1> */ input  pag4_page_ok_l,
  /* <dl1> */ input  pag4_page_refill_l,
  /* <ed2> */ input  phase_change_coming_l,
  /* <fp2> */ input  pma5_csh_writeback_cyc_l,
  /* <bm2> */ input  pma5_page_refill_cyc_l,
  /* <de1> */ input  vma1_ac_ref_a_h
);

`include "csh23nets.svh"

endmodule	// csh23
