module tapped_delay_50_10(input bit in, output bit t1,t2,t3,t4, out);
  always_comb t1 = in;
  always_comb t2 = in;
  always_comb t3 = in;
  always_comb t4 = in;
  always_comb out = in;
endmodule // tapped_delay_50_10
