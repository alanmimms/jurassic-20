module chx;
`include "chx.svh"
endmodule	// chx
