module zero6(output bit q1, q2, q3, q4, q5, q6);
  always_comb begin
    q1 = 0;
    q2 = 0;
    q3 = 0;
    q4 = 0;
    q5 = 0;
    q6 = 0;
  end
endmodule // just_six_zero
