module shm;
`include "shm.svh"
endmodule	// shm
