module mb015(
      input  ar_06_a_h                         /* <fc1> */,
      input  ar_07_a_h                         /* <fd1> */,
      input  ar_08_a_h                         /* <eu2> */,
      input  ar_09_a_h                         /* <ev2> */,
      input  ar_10_a_h                         /* <cv2> */,
      input  ar_11_a_h                         /* <bu2> */,
      input  ar_24_a_h                         /* <dd2> */,
      input  ar_25_a_h                         /* <cs2> */,
      input  ar_26_a_h                         /* <bp1> */,
      input  ar_27_a_h                         /* <bj2> */,
      input  ar_28_a_h                         /* <bm2> */,
      input  ar_29_a_h                         /* <bf1> */,
      input  cache_data_06_a_h                 /* <er2> */,
      input  cache_data_07_a_h                 /* <ef1> */,
      input  cache_data_08_a_h                 /* <ff2> */,
      input  cache_data_09_a_h                 /* <er1> */,
      input  cache_data_10_a_h                 /* <cr1> */,
      input  cache_data_11_a_h                 /* <cm2> */,
      input  cache_data_24_a_h                 /* <dk2> */,
      input  cache_data_25_a_h                 /* <dk1> */,
      input  cache_data_26_a_h                 /* <am1> */,
      input  cache_data_27_a_h                 /* <ak1> */,
      input  cache_data_28_a_h                 /* <ar1> */,
      input  cache_data_29_a_h                 /* <ap1> */,
      input  cbus_d06_re_h                     /* <cj1> */,
      output cbus_d06_te_h                     /* <ee1> */,
      input  cbus_d07_re_h                     /* <cj2> */,
      output cbus_d07_te_h                     /* <ee2> */,
      input  cbus_d08_re_h                     /* <bs2> */,
      output cbus_d08_te_h                     /* <el2> */,
      input  cbus_d09_re_h                     /* <bc1> */,
      output cbus_d09_te_h                     /* <em1> */,
      input  cbus_d10_re_h                     /* <br1> */,
      output cbus_d10_te_h                     /* <df1> */,
      input  cbus_d11_re_h                     /* <bd2> */,
      output cbus_d11_te_h                     /* <dl2> */,
      input  cbus_d24_re_h                     /* <ch2> */,
      output cbus_d24_te_h                     /* <dn1> */,
      input  cbus_d25_re_h                     /* <cf1> */,
      output cbus_d25_te_h                     /* <dm2> */,
      input  cbus_d26_re_h                     /* <be2> */,
      output cbus_d26_te_h                     /* <ah2> */,
      input  cbus_d27_re_h                     /* <bj1> */,
      output cbus_d27_te_h                     /* <af2> */,
      input  cbus_d28_re_h                     /* <be1> */,
      output cbus_d28_te_h                     /* <aj2> */,
      input  cbus_d29_re_h                     /* <bl1> */,
      output cbus_d29_te_h                     /* <ak2> */,
      input  ccl_ccw_buf_wr_l                  /* <fk1> */,
      input  ccl_ch_buf_en_l                   /* <ae2> */,
      input  ccl_mix_mb_sel_h                  /* <es1> */,
      input  ccw_buf_06_in_h                   /* <fl1> */,
      input  ccw_buf_07_in_h                   /* <fm2> */,
      input  ccw_buf_08_in_h                   /* <fh2> */,
      input  ccw_buf_09_in_h                   /* <fj2> */,
      input  ccw_buf_10_in_h                   /* <cl2> */,
      input  ccw_buf_11_in_h                   /* <cl1> */,
      input  ccw_buf_24_in_h                   /* <ck2> */,
      input  ccw_buf_25_in_h                   /* <ck1> */,
      input  ccw_buf_26_in_h                   /* <at2> */,
      input  ccw_buf_27_in_h                   /* <as1> */,
      input  ccw_buf_28_in_h                   /* <ap2> */,
      input  ccw_buf_29_in_h                   /* <am2> */,
      input  ccw_buf_adr_0_h                   /* <fk2> */,
      input  ccw_buf_adr_1_h                   /* <fj1> */,
      input  ccw_buf_adr_2_h                   /* <fl2> */,
      input  ccw_buf_adr_3_h                   /* <fm1> */,
      output ccw_mix_06_h                      /* <ek2> */,
      output ccw_mix_07_h                      /* <eh2> */,
      output ccw_mix_08_h                      /* <ff1> */,
      output ccw_mix_09_h                      /* <es2> */,
      output ccw_mix_10_h                      /* <cp2> */,
      output ccw_mix_11_h                      /* <cn1> */,
      output ccw_mix_24_h                      /* <dl1> */,
      output ccw_mix_25_h                      /* <dh2> */,
      output ccw_mix_26_h                      /* <al2> */,
      output ccw_mix_27_h                      /* <al1> */,
      output ccw_mix_28_h                      /* <as2> */,
      output ccw_mix_29_h                      /* <ar2> */,
      input  ch_buf_wr_04_l                    /* <aj1> */,
      input  ch_buf_wr_1_l                     /* <ep1> */,
      input  ch_reverse_h                      /* <bd1> */,
      input  ch_t0_l                           /* <fs2> */,
      input  ch_t2_l                           /* <af1> */,
      input  clk_mb_06_h                       /* <cr2> */,
      input  con_ki10_paging_mode_l            /* <ek1> */,
      input  crc_buf_mb_sel_h                  /* <dt2> */,
      input  crc_cbus_out_hold_h               /* <fu2> */,
      input  crc_ch_buf_adr_0_h                /* <fp2> */,
      input  crc_ch_buf_adr_1_h                /* <fr2> */,
      input  crc_ch_buf_adr_2_h                /* <fp1> */,
      input  crc_ch_buf_adr_3_h                /* <de1> */,
      input  crc_ch_buf_adr_4_h                /* <dj1> */,
      input  crc_ch_buf_adr_5_h                /* <de2> */,
      input  crc_ch_buf_adr_6_h                /* <ae1> */,
      input  mb0_hold_in_h                     /* <ad2> */,
      input  mb1_hold_in_h                     /* <ad1> */,
      input  mb2_hold_in_h                     /* <aa1> */,
      input  mb3_hold_in_h                     /* <ac1> */,
      output mb_06_h                           /* <fd2> */,
      output mb_06to11_par_odd_h               /* <ds2> */,
      output mb_07_h                           /* <dr2> */,
      output mb_08_h                           /* <dp2> */,
      output mb_09_h                           /* <dm1> */,
      output mb_10_h                           /* <dr1> */,
      output mb_11_h                           /* <dp1> */,
      output mb_24_h                           /* <av2> */,
      output mb_24to29_par_odd_h               /* <au2> */,
      output mb_25_h                           /* <ba1> */,
      output mb_26_h                           /* <cd2> */,
      output mb_27_h                           /* <cd1> */,
      output mb_28_h                           /* <ca1> */,
      output mb_29_h                           /* <bv2> */,
      input  mb_in_sel_1_h                     /* <ej1> */,
      input  mb_in_sel_2_h                     /* <el1> */,
      input  mb_in_sel_4_h                     /* <ep2> */,
      input  mb_sel_1_en_h                     /* <fr1> */,
      input  mb_sel_2_en_h                     /* <ft2> */,
      input  mb_sel_hold_h                     /* <fv2> */,
      input  mem_data_in_06_h                  /* <em2> */,
      input  mem_data_in_07_h                  /* <ej2> */,
      input  mem_data_in_08_h                  /* <ea1> */,
      input  mem_data_in_09_h                  /* <dv2> */,
      input  mem_data_in_10_h                  /* <cp1> */,
      input  mem_data_in_11_h                  /* <cm1> */,
      input  mem_data_in_24_h                  /* <dj2> */,
      input  mem_data_in_25_h                  /* <df2> */,
      input  mem_data_in_26_h                  /* <bm1> */,
      input  mem_data_in_27_h                  /* <bk2> */,
      input  mem_data_in_28_h                  /* <bl2> */,
      input  mem_data_in_29_h                  /* <bk1> */,
      input  mem_to_c_en_l                     /* <ed2> */,
      input  mem_to_c_sel_1_h                  /* <ed1> */,
      input  mem_to_c_sel_2_h                  /* <ds1> */,
      output mem_to_cache_06_h                 /* <en1> */,
      output mem_to_cache_07_h                 /* <ef2> */,
      output mem_to_cache_08_h                 /* <ec1> */,
      output mem_to_cache_09_h                 /* <du2> */,
      output mem_to_cache_10_h                 /* <cf2> */,
      output mem_to_cache_11_h                 /* <cc1> */,
      output mem_to_cache_24_h                 /* <cs1> */,
      output mem_to_cache_25_h                 /* <dd1> */,
      output mem_to_cache_26_h                 /* <br2> */,
      output mem_to_cache_27_h                 /* <bf2> */,
      output mem_to_cache_28_h                 /* <bp2> */,
      output mem_to_cache_29_h                 /* <bh2> */,
      input  nxm_any_l                         /* <fs1> */,
      output pt_in_06_h                        /* <fe1> */,
      output pt_in_07_h                        /* <fe2> */,
      output pt_in_08_h                        /* <fa1> */,
      output pt_in_09_h                        /* <et2> */,
      output pt_in_10_h                        /* <dc1> */,
      output pt_in_11_h                        /* <da1> */,
      output pt_in_24_h                        /* <cu2> */,
      output pt_in_25_h                        /* <ct2> */,
      output pt_in_26_h                        /* <ce1> */,
      output pt_in_27_h                        /* <ce2> */,
      output pt_in_28_h                        /* <bs1> */,
      output pt_in_29_h                        /* <bt2> */
);

`include "mb015nets.svh"

endmodule	// mb015
