module pma;
`include "pma.svh"
endmodule	// pma
