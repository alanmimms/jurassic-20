module apr;
`include "apr.svh"
endmodule	// apr
