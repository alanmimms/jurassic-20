module edp51(
  /* <cp2> */ input  ad_04_h,
  /* <el2> */ input  ad_05_h,
  /* <ck1> */ output ad_06_a_h,
  /* <cn1> */ output ad_06_a_l,
  /* <ep2> */ output ad_06_h,
  /* <at2> */ output ad_06to11Eq0_l,
  /* <dl1> */ output ad_07_h,
  /* <dr2> */ output ad_08_h,
  /* <dr1> */ output ad_09_h,
  /* <cf2> */ output ad_10_a_h,
  /* <cp1> */ output ad_10_h,
  /* <ce1> */ output ad_11_a_h,
  /* <el1> */ output ad_11_h,
  /* <ep1> */ input  ad_12_h,
  /* <am1> */ output ad_cg_06_h,
  /* <am2> */ output ad_cg_08_h,
  /* <aj1> */ output ad_cp_06_h,
  /* <af1> */ output ad_cp_08_h,
  /* <cu2> */ output ad_cry_07_h,
  /* <ct2> */ output ad_cry_07_l,
  /* <al1> */ input  ad_cry_12_h,
  /* <cv2> */ output ad_ex_04_h,
  /* <cr1> */ output ad_ex_05_h,
  /* <cl2> */ output ad_overflow_06_l,
  /* <es2> */ input  adx_05_h,
  /* <cf1> */ output adx_06_a_h,
  /* <cj2> */ output adx_06_h,
  /* <dk1> */ output adx_10_h,
  /* <es1> */ output adx_11_h,
  /* <cj1> */ input  adx_12_h,
  /* <al2> */ output adx_cg_06_h,
  /* <ak2> */ output adx_cg_09_h,
  /* <ae1> */ output adx_cp_06_h,
  /* <af2> */ output adx_cp_09_h,
  /* <ak1> */ input  adx_cry_12_h,
  /* <fr2> */ input  apr_fm_adr_10_h,
  /* <fp2> */ input  apr_fm_adr_1_h,
  /* <fs1> */ input  apr_fm_adr_2_h,
  /* <fn1> */ input  apr_fm_adr_4_h,
  /* <fr1> */ input  apr_fm_block_1_h,
  /* <fm1> */ input  apr_fm_block_2_h,
  /* <fp1> */ input  apr_fm_block_4_h,
  /* <fj2> */ output ar_06_a_h,
  /* <ft2> */ output ar_06_b_h,
  /* <fs2> */ output ar_06_c_h,
  /* <dm2> */ output ar_06_d_h,
  /* <bk2> */ output ar_06_h,
  /* <fc1> */ output ar_07_a_h,
  /* <fu2> */ output ar_07_b_h,
  /* <fv2> */ output ar_07_c_h,
  /* <bl2> */ output ar_07_h,
  /* <ff2> */ output ar_08_a_h,
  /* <cl1> */ output ar_08_b_h,
  /* <ch2> */ output ar_08_c_h,
  /* <eu2> */ output ar_09_a_h,
  /* <ck2> */ output ar_09_b_h,
  /* <cm1> */ output ar_09_c_h,
  /* <ev2> */ output ar_10_a_h,
  /* <fk1> */ output ar_10_b_h,
  /* <fk2> */ output ar_10_c_h,
  /* <et2> */ output ar_11_a_h,
  /* <fl2> */ output ar_11_b_h,
  /* <fl1> */ output ar_11_c_h,
  /* <bk1> */ input  ar_12_h,
  /* <bl1> */ input  ar_13_h,
  /* <em2> */ input  armm_06_h,
  /* <ea1> */ input  armm_07_h,
  /* <ee1> */ input  armm_08_h,
  /* <dd2> */ input  armm_09_h,
  /* <de1> */ input  armm_10_h,
  /* <ef2> */ input  armm_11_h,
  /* <as2> */ output arx_06_a_h,
  /* <br2> */ output arx_06_b_h,
  /* <ej2> */ output arx_06_h,
  /* <as1> */ output arx_07_a_h,
  /* <cm2> */ output arx_07_b_h,
  /* <bd2> */ output arx_07_h,
  /* <dc1> */ output arx_08_h,
  /* <aj2> */ output arx_09_h,
  /* <ac1> */ output arx_10_h,
  /* <aa1> */ output arx_11_h,
  /* <ej1> */ input  arx_12_h,
  /* <bd1> */ input  arx_13_h,
  /* <bm2> */ output br_06_a_h,
  /* <bm1> */ input  br_12_a_h,
  /* <be2> */ output brx_06_h,
  /* <be1> */ input  brx_12_h,
  /* <em1> */ input  cache_data_06_b_h,
  /* <ed2> */ input  cache_data_07_b_h,
  /* <ee2> */ input  cache_data_08_b_h,
  /* <dd1> */ input  cache_data_09_b_h,
  /* <dl2> */ input  cache_data_10_b_h,
  /* <cc1> */ input  cache_data_11_b_h,
  /* <cr2> */ input  clk_edp_06_h,
  /* <ce2> */ input  con_fm_write_00to17_l,
  /* <ar1> */ input  cram_Nr_06_h,
  /* <ap1> */ input  cram_Nr_07_h,
  /* <ba1> */ input  cram_Nr_08_h,
  /* <ap2> */ input  cram_Nr_09_h,
  /* <av2> */ input  cram_Nr_10_h,
  /* <au2> */ input  cram_Nr_11_h,
  /* <an1> */ input  cram_ad_boole_06_h,
  /* <ad2> */ input  cram_ad_sel_1_06_h,
  /* <ah2> */ input  cram_ad_sel_2_06_h,
  /* <ae2> */ input  cram_ad_sel_4_06_h,
  /* <ad1> */ input  cram_ad_sel_8_06_h,
  /* <bn1> */ input  cram_ada_dis_06_h,
  /* <bj1> */ input  cram_ada_sel_1_06_h,
  /* <bf2> */ input  cram_ada_sel_2_06_h,
  /* <bt2> */ input  cram_adb_sel_1_06_h,
  /* <bt1> */ input  cram_adb_sel_1_06_h,
  /* <bs1> */ input  cram_adb_sel_2_06_h,
  /* <ff1> */ input  cram_arxm_sel_4_00_h,
  /* <dj2> */ input  cram_br_load_a_h,
  /* <ar2> */ input  cram_brx_load_a_h,
  /* <fe2> */ input  ctl_ad_to_ebus_l_h,
  /* <dh2> */ input  ctl_ar_00to08_load_l,
  /* <eh2> */ input  ctl_ar_00to11_clr_h,
  /* <ek2> */ input  ctl_ar_09to17_load_l,
  /* <en1> */ input  ctl_arl_sel_1_h,
  /* <ek1> */ input  ctl_arl_sel_2_h,
  /* <er1> */ input  ctl_arl_sel_4_h,
  /* <br1> */ input  ctl_arx_load_h,
  /* <fj1> */ input  ctl_arxl_sel_1_h,
  /* <fd2> */ input  ctl_arxl_sel_2_h,
  /* <bu2> */ input  ctl_mq_sel_1_h,
  /* <bv2> */ input  ctl_mq_sel_2_h,
  /* <dn1> */ input  ctl_mqm_en_h,
  /* <dj1> */ input  ctl_mqm_sel_1_h,
  /* <dm1> */ input  ctl_mqm_sel_2_h,
  /* <fd1> */ input  diag_04_a_h,
  /* <fa1> */ input  diag_05_a_h,
  /* <fe1> */ input  diag_06_a_h,
  /* <ef1> */ input  diag_read_func_12x_h,
  /* <dv2> */ output ebus_d06_e_h,
  /* <ds2> */ output ebus_d07_e_h,
  /* <dt2> */ output ebus_d08_e_h,
  /* <dp1> */ output ebus_d09_e_h,
  /* <dp2> */ output ebus_d10_e_h,
  /* <du2> */ output ebus_d11_e_h,
  /* <fm2> */ output edp_fm_parity_06to11_h,
  /* <cs2> */ input  mq_04_h,
  /* <cd2> */ output mq_06_h,
  /* <cs1> */ output mq_10_h,
  /* <df1> */ output mq_11_h,
  /* <cd1> */ input  mq_12_h,
  /* <ed1> */ input  sh_06_h,
  /* <ec1> */ input  sh_07_h,
  /* <ds1> */ input  sh_08_h,
  /* <da1> */ input  sh_09_h,
  /* <de2> */ input  sh_10_h,
  /* <ca1> */ input  sh_11_h,
  /* <bj2> */ input  vma_held_or_pc_06_h,
  /* <bh2> */ input  vma_held_or_pc_07_h,
  /* <bf1> */ input  vma_held_or_pc_08_h,
  /* <bp2> */ input  vma_held_or_pc_09_h,
  /* <bp1> */ input  vma_held_or_pc_10_h,
  /* <bc1> */ input  vma_held_or_pc_11_h
);

`include "edp51nets.svh"

endmodule	// edp51
