module mbz20(
  /* <fv2> */  input a_change_coming_in_l,
  /* <ep2> */  input ackn_pulse_l,
  /* <fe1> */  input apr_any_ebox_err_flg_h,
  /* <al2> */  input apr_ebox_era_h,
  /* <eu2> */  input apr_ebox_sbus_diag_l,
  /* <au2> */  input apr_mb_par_err_l,
  /* <dl1> */  input apr_nxm_err_l,
  /* <at2> */  input apr_sbus_err_l,
  /* <br1> */  input cache_to_mb_t4_l,
  /* <dk1> */  input cbus_par_left_re_h,
  /* <ce1> */ output cbus_par_left_te_h,
  /* <dj2> */  input cbus_par_right_re_h,
  /* <cd1> */ output cbus_par_right_te_h,
  /* <da1> */  input ccl_ch_test_mb_par_l,
  /* <dt2> */  input ccl_chan_ept_h,
  /* <bh2> */  input ccl_chan_to_mem_l,
  /* <dj1> */  input ccl_data_reverse_h,
  /* <dc1> */  input ccl_hold_mem_h,
  /* <es1> */  input ccl_odd_wc_par_h,
  /* <et2> */  input ccw_odd_adr_par_h,
  /* <ek2> */  input ch_buf_wr_06_l,
  /* <ft2> */  input ch_t0_l,
  /* <ek1> */  input ch_t2_l,
  /* <cj1> */ output chan_adr_par_err_l,
  /* <fk1> */ output chan_nxm_err_l,
  /* <cf2> */ output chan_par_err_l,
  /* <cm2> */ output chan_read_h,
  /* <cu2> */ output chan_read_l,
  /* <cr2> */  input clk_mbz_h,
  /* <ea1> */  input core_busy_a_h,
  /* <dm2> */ output core_busy_h,
  /* <dh2> */ output core_busy_l,
  /* <ef1> */  input core_rd_in_prog_h,
  /* <fr2> */  input crc_buf_mb_sel_h,
  /* <cc1> */  input crc_cbus_out_hold_h,
  /* <ej1> */  input crc_ch_buf_adr_0_h,
  /* <ef2> */  input crc_ch_buf_adr_1_h,
  /* <eh2> */  input crc_ch_buf_adr_2_h,
  /* <fs2> */  input crc_ch_buf_adr_3_h,
  /* <ee1> */  input crc_ch_buf_adr_4_h,
  /* <ee2> */  input crc_ch_buf_adr_5_h,
  /* <em2> */  input crc_ch_buf_adr_6_h,
  /* <ds2> */  input csh_chan_cyc_l,
  /* <ej2> */  input csh_ebox_cyc_a_l,
  /* <es2> */ output csh_en_csh_data_l,
  /* <fe2> */  input csh_par_bit_00_a_h,
  /* <fc1> */  input csh_par_bit_00_b_h,
  /* <fh2> */  input csh_par_bit_01_a_h,
  /* <fd1> */  input csh_par_bit_01_b_h,
  /* <ff1> */  input csh_par_bit_02_a_h,
  /* <fj2> */  input csh_par_bit_02_b_h,
  /* <ff2> */  input csh_par_bit_03_a_h,
  /* <fd2> */  input csh_par_bit_03_b_h,
  /* <fs1> */ output csh_par_bit_a_h,
  /* <fa1> */ output csh_par_bit_b_h,
  /* <ct2> */ output csh_par_bit_in_h,
  /* <ah2> */  input diag_05_b_h,
  /* <af2> */  input diag_06_b_h,
  /* <fm1> */  input diag_load_func_071_l,
  /* <dr2> */  input diag_read_func_16x_l,
  /* <er1> */  input e_cache_wr_cyc_l,
  /* <bu2> */ output ebus_d00_e_h,
  /* <bv2> */ output ebus_d01_e_h,
  /* <bs1> */ output ebus_d02_e_h,
  /* <bp1> */ output ebus_d03_e_h,
  /* <ca1> */ output ebus_d04_e_h,
  /* <bt2> */ output ebus_d05_e_h,
  /* <bp2> */ output ebus_d06_e_h,
  /* <bn1> */ output ebus_d07_e_h,
  /* <ch2> */ output ebus_d08_e_h,
  /* <cl1> */ output ebus_d14_e_h,
  /* <cj2> */ output ebus_d15_e_h,
  /* <cd2> */ output ebus_d16_e_h,
  /* <cp1> */ output ebus_d17_e_h,
  /* <cn1> */ output ebus_d18_e_h,
  /* <cp2> */ output ebus_d19_e_h,
  /* <cl2> */ output ebus_d20_e_h,
  /* <df1> */ output ebus_d21_e_h,
  /* <dl2> */ output ebus_d22_e_h,
  /* <df2> */ output ebus_d23_e_h,
  /* <dd2> */ output ebus_d24_e_h,
  /* <ec1> */ output ebus_d25_e_h,
  /* <dm1> */ output ebus_d26_e_h,
  /* <fp1> */ output ebus_d34_e_h,
  /* <ce2> */ output ebus_d35_e_h,
  /* <fk2> */ output hi,
  /* <aa1> */ output hold_era_h,
  /* <ad1> */  input load_ebus_reg_l,
  /* <ad2> */  input mb_data_code_1_h,
  /* <af1> */  input mb_data_code_2_h,
  /* <ep1> */ output mb_in_sel_1_h,
  /* <fu2> */ output mb_in_sel_2_h,
  /* <er2> */ output mb_in_sel_4_h,
  /* <cm1> */ output mb_par_bit_in_h,
  /* <en1> */  input mb_par_h,
  /* <av2> */  input mb_par_odd_h,
  /* <ar1> */  input mb_req_hold_h,
  /* <ae1> */  input mb_sel_1_h,
  /* <ae2> */  input mb_sel_2_h,
  /* <ac1> */  input mb_test_par_a_in_l,
  /* <fr1> */ output mbox_adr_par_err_l,
  /* <bm2> */ output mbox_mb_par_err_l,
  /* <fp2> */ output mbox_nxm_err_l,
  /* <de1> */ output mbox_sbus_err_l,
  /* <ds1> */ output mbz1_rdNgpseNgwr_ref_l,
  /* <bm1> */  input mcl_vma_user_h,
  /* <ar2> */  input mem_adr_par_err_h,
  /* <du2> */ output mem_busy_h,
  /* <ap2> */  input mem_error_h,
  /* <cs2> */  input mem_par_in_h,
  /* <aj2> */  input mem_rd_rq_b_h,
  /* <fl2> */  input mem_start_a_h,
  /* <fm2> */  input mem_start_b_h,
  /* <cv2> */ output mem_to_c_diag_en_l,
  /* <el2> */  input mem_to_c_en_l,
  /* <fj1> */  input mem_to_c_sel_1_h,
  /* <el1> */  input mem_to_c_sel_2_h,
  /* <br2> */  input mem_wr_rq_l,
  /* <dn1> */  input mr_reset_06_h,
  /* <ed2> */  input mtr_cca_writeback_l,
  /* <ck2> */ output nxm_ackn_h,
  /* <de2> */ output nxm_any_l,
  /* <dr1> */ output nxm_data_val_l,
  /* <dp1> */  input pag_mb_00to17_par_h,
  /* <dp2> */  input pag_mb_18to35_par_h,
  /* <bf2> */  input paged_ref_h,
  /* <bl2> */  input pf_hold_01_in_h,
  /* <bl1> */  input pf_hold_02_in_h,
  /* <bk1> */  input pf_hold_03_in_h,
  /* <bf1> */  input pf_hold_04_in_h,
  /* <as1> */  input pf_hold_05_in_h,
  /* <bs2> */  input phase_change_coming_l,
  /* <bn2> */  input pma_14_h,
  /* <bj1> */  input pma_15_h,
  /* <bk2> */  input pma_16_h,
  /* <bd2> */  input pma_17_h,
  /* <bc1> */  input pma_18_h,
  /* <ba1> */  input pma_19_h,
  /* <bd1> */  input pma_20_h,
  /* <am1> */  input pma_21_h,
  /* <am2> */  input pma_22_h,
  /* <an1> */  input pma_23_h,
  /* <as2> */  input pma_24_h,
  /* <al1> */  input pma_25_h,
  /* <ak1> */  input pma_26_h,
  /* <ak2> */  input pma_34_h,
  /* <ap1> */  input pma_35_h,
  /* <be1> */  input pt_cache_h,
  /* <be2> */  input pt_public_h,
  /* <fn1> */  input rq_hold_ff_h,
  /* <cr1> */  input sh_ar_par_odd_a_h
);

`include "mbz20nets.svh"

endmodule	// mbz20
