module crc;
`include "crc.svh"
endmodule	// crc
