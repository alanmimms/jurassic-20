module mbc;
`include "mbc.svh"
endmodule	// mbc
