module mcl;
`include "mcl.svh"
endmodule	// mcl
