module tapped_delay_50_10(input bit in, output bit t1,t2,t3,t4, out);
  assign t1 = in;
  assign t2 = in;
  assign t3 = in;
  assign t4 = in;
  assign out = in;
endmodule // tapped_delay_50_10
