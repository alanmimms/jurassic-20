module edp53(
      output ad_00_a_h                         /* <ck1> */,
      output ad_00_a_l                         /* <cn1> */,
      output ad_00_h                           /* <ep2> */,
      output ad_00to05Eq0_l                    /* <at2> */,
      output ad_01_h                           /* <dl1> */,
      output ad_02_h                           /* <dr2> */,
      output ad_03_h                           /* <dr1> */,
      output ad_04_a_h                         /* <cf2> */,
      output ad_04_h                           /* <cp1> */,
      output ad_05_a_h                         /* <ce1> */,
      output ad_05_h                           /* <el1> */,
      input  ad_06_h                           /* <ep1> */,
      input  ad_35_h                           /* <es2> */,
      output ad_cg_00_h                        /* <am1> */,
      output ad_cg_02_h                        /* <am2> */,
      output ad_cp_00_h                        /* <aj1> */,
      output ad_cp_02_h                        /* <af1> */,
      output ad_cry_01_h                       /* <cu2> */,
      output ad_cry_01_l                       /* <ct2> */,
      input  ad_cry_06_h                       /* <al1> */,
      input  ad_ex_Ng01_h                      /* <el2><cr1> */,
      input  ad_ex_Ng02_h                      /* <cp2><cv2> */,
      output ad_overflow_00_l                  /* <cl2> */,
      output adx_00_a_h                        /* <cf1> */,
      output adx_00_h                          /* <cj2> */,
      output adx_04_h                          /* <dk1> */,
      output adx_05_h                          /* <es1> */,
      input  adx_06_h                          /* <cj1> */,
      input  adx_34_h                          /* <cs2> */,
      output adx_cg_00_h                       /* <al2> */,
      output adx_cg_03_h                       /* <ak2> */,
      output adx_cp_00_h                       /* <ae1> */,
      output adx_cp_03_h                       /* <af2> */,
      input  adx_cry_06_h                      /* <ak1> */,
      input  apr_fm_adr_10_h                   /* <fr2> */,
      input  apr_fm_adr_1_h                    /* <fp2> */,
      input  apr_fm_adr_2_h                    /* <fs1> */,
      input  apr_fm_adr_4_h                    /* <fn1> */,
      input  apr_fm_block_1_h                  /* <fr1> */,
      input  apr_fm_block_2_h                  /* <fm1> */,
      input  apr_fm_block_4_h                  /* <fp1> */,
      output ar_00_a_h                         /* <fj2> */,
      output ar_00_b_h                         /* <ft2> */,
      output ar_00_c_h                         /* <fs2> */,
      output ar_00_d_h                         /* <dm2> */,
      output ar_00_h                           /* <bk2> */,
      output ar_01_a_h                         /* <fc1> */,
      output ar_01_b_h                         /* <fu2> */,
      output ar_01_c_h                         /* <fv2> */,
      output ar_01_h                           /* <bl2> */,
      output ar_02_a_h                         /* <ff2> */,
      output ar_02_b_h                         /* <cl1> */,
      output ar_02_c_h                         /* <ch2> */,
      output ar_03_a_h                         /* <eu2> */,
      output ar_03_b_h                         /* <ck2> */,
      output ar_03_c_h                         /* <cm1> */,
      output ar_04_a_h                         /* <ev2> */,
      output ar_04_b_h                         /* <fk1> */,
      output ar_04_c_h                         /* <fk2> */,
      output ar_05_a_h                         /* <et2> */,
      output ar_05_b_h                         /* <fl2> */,
      output ar_05_c_h                         /* <fl1> */,
      input  ar_06_h                           /* <bk1> */,
      input  ar_07_h                           /* <bl1> */,
      input  armm_00_h                         /* <em2> */,
      input  armm_01_h                         /* <ea1> */,
      input  armm_02_h                         /* <ee1> */,
      input  armm_03_h                         /* <dd2> */,
      input  armm_04_h                         /* <de1> */,
      input  armm_05_h                         /* <ef2> */,
      output arx_00_a_h                        /* <as2> */,
      output arx_00_b_h                        /* <br2> */,
      output arx_00_h                          /* <ej2> */,
      output arx_01_a_h                        /* <as1> */,
      output arx_01_b_h                        /* <cm2> */,
      output arx_01_h                          /* <bd2> */,
      output arx_02_h                          /* <dc1> */,
      output arx_03_h                          /* <aj2> */,
      output arx_04_h                          /* <ac1> */,
      output arx_05_h                          /* <aa1> */,
      input  arx_06_h                          /* <ej1> */,
      input  arx_07_h                          /* <bd1> */,
      output br_00_a_h                         /* <bm2> */,
      input  br_06_a_h                         /* <bm1> */,
      output brx_00_h                          /* <be2> */,
      input  brx_06_h                          /* <be1> */,
      input  cache_data_00_b_h                 /* <em1> */,
      input  cache_data_01_b_h                 /* <ed2> */,
      input  cache_data_02_b_h                 /* <ee2> */,
      input  cache_data_03_b_h                 /* <dd1> */,
      input  cache_data_04_b_h                 /* <dl2> */,
      input  cache_data_05_b_h                 /* <cc1> */,
      input  clk_edp_00_h                      /* <cr2> */,
      input  con_fm_write_00to17_l             /* <ce2> */,
      input  cram_Nr_00_h                      /* <ar1> */,
      input  cram_Nr_01_h                      /* <ap1> */,
      input  cram_Nr_02_h                      /* <ba1> */,
      input  cram_Nr_03_h                      /* <ap2> */,
      input  cram_Nr_04_h                      /* <av2> */,
      input  cram_Nr_05_h                      /* <au2> */,
      input  cram_ad_boole_00_h                /* <an1> */,
      input  cram_ad_sel_1_00_h                /* <ad2> */,
      input  cram_ad_sel_2_00_h                /* <ah2> */,
      input  cram_ad_sel_4_00_h                /* <ae2> */,
      input  cram_ad_sel_8_00_h                /* <ad1> */,
      input  cram_ada_dis_00_h                 /* <bn1> */,
      input  cram_ada_sel_1_00_h               /* <bj1> */,
      input  cram_ada_sel_2_00_h               /* <bf2> */,
      input  cram_adb_sel_1_00_h               /* <bt2> */,
      input  cram_adb_sel_2_00_h               /* <bs1> */,
      input  cram_arxm_sel_4_00_h              /* <ff1> */,
      input  cram_br_load_a_h                  /* <dj2> */,
      input  cram_brx_load_a_h                 /* <ar2> */,
      input  ctl_ad_to_ebus_l_h                /* <fe2> */,
      input  ctl_ar_00to08_load_l              /* <ek2><dh2> */,
      input  ctl_ar_00to11_clr_h               /* <eh2> */,
      input  ctl_arl_sel_1_h                   /* <en1> */,
      input  ctl_arl_sel_2_h                   /* <ek1> */,
      input  ctl_arl_sel_4_h                   /* <er1> */,
      input  ctl_arx_load_h                    /* <br1> */,
      input  ctl_arxl_sel_1_h                  /* <fj1> */,
      input  ctl_arxl_sel_2_h                  /* <fd2> */,
      input  ctl_mq_sel_1_h                    /* <bu2> */,
      input  ctl_mq_sel_2_h                    /* <bv2> */,
      input  ctl_mqm_en_h                      /* <dn1> */,
      input  ctl_mqm_sel_1_h                   /* <dj1> */,
      input  ctl_mqm_sel_2_h                   /* <dm1> */,
      input  diag_04_a_h                       /* <fd1> */,
      input  diag_05_a_h                       /* <fa1> */,
      input  diag_06_a_h                       /* <fe1> */,
      input  diag_read_func_12x_h              /* <ef1> */,
      output ebus_d00_e_h                      /* <dv2> */,
      output ebus_d01_e_h                      /* <ds2> */,
      output ebus_d02_e_h                      /* <dt2> */,
      output ebus_d03_e_h                      /* <dp1> */,
      output ebus_d04_e_h                      /* <dp2> */,
      output ebus_d05_e_h                      /* <du2> */,
      output edp_fm_parity_00to05_h            /* <fm2> */,
      input  hi                                /* <bs2> */,
      output mq_00_h                           /* <cd2> */,
      output mq_04_h                           /* <cs1> */,
      output mq_05_h                           /* <df1> */,
      input  mq_06_h                           /* <cd1> */,
      input  sh_00_h                           /* <ed1> */,
      input  sh_01_h                           /* <ec1> */,
      input  sh_02_h                           /* <ds1> */,
      input  sh_03_h                           /* <da1> */,
      input  sh_04_h                           /* <de2> */,
      input  sh_05_h                           /* <ca1> */,
      input  vma_held_or_pc_00_h               /* <bj2> */,
      input  vma_held_or_pc_01_h               /* <bh2> */,
      input  vma_held_or_pc_02_h               /* <bf1> */,
      input  vma_held_or_pc_03_h               /* <bp2> */,
      input  vma_held_or_pc_04_h               /* <bp1> */,
      input  vma_held_or_pc_05_h               /* <bc1> */
);

`include "edp53nets.svh"

endmodule	// edp53
