module ccl11(
      output ccl_act_flag_clr_l                /* <be2> */,
      output ccl_act_flag_req_l                /* <bd1> */,
      output ccl_af_wd0_req_h                  /* <fc1> */,
      output ccl_af_wd1_req_h                  /* <fa1> */,
      output ccl_af_wd2_req_h                  /* <fh2> */,
      output ccl_af_wd3_req_h                  /* <fj2> */,
      output ccl_alu_minus_l                   /* <ee1> */,
      output ccl_alu_plus_l                    /* <aj2> */,
      output ccl_buf_adr_3_h                   /* <ej1> */,
      output ccl_ccw_buf_wr_l                  /* <bt2> */,
      output ccl_ccw_reg_load_h                /* <cu2> */,
      output ccl_ccwf_clr_h                    /* <aj1> */,
      output ccl_ccwf_clr_l                    /* <av2> */,
      output ccl_ccwf_req_h                    /* <ek2> */,
      output ccl_ch_buf_wr_en_l                /* <bs2> */,
      output ccl_ch_load_mb_l                  /* <dk2> */,
      output ccl_ch_mb_sel_1_h                 /* <ee2> */,
      output ccl_ch_mb_sel_2_h                 /* <ds2> */,
      output ccl_ch_test_mb_par_l              /* <dl2> */,
      output ccl_chan_ept_h                    /* <eh2> */,
      output ccl_chan_ept_l                    /* <ar1> */,
      output ccl_chan_req_h                    /* <dv2> */,
      output ccl_chan_req_l                    /* <df2> */,
      output ccl_chan_to_mem_h                 /* <dd1> */,
      output ccl_chan_to_mem_l                 /* <df1> */,
      output ccl_cons_0_h                      /* <fv2> */,
      output ccl_cons_1_h                      /* <ft2> */,
      output ccl_cons_2_h                      /* <fu2> */,
      output ccl_csh_chan_cyc_h                /* <ef1> */,
      output ccl_data_reverse_h                /* <cp2> */,
      output ccl_err_req_l                     /* <ae2> */,
      output ccl_error_h                       /* <ba1> */,
      output ccl_hold_mem_h                    /* <bs1> */,
      output ccl_last_xfer_err_in_h            /* <er2> */,
      output ccl_load_ac_h                     /* <ct2> */,
      output ccl_load_ac_l                     /* <cs2> */,
      output ccl_mb_cyc_t2_l                   /* <el1> */,
      output ccl_mb_req_t2_l                   /* <ek1> */,
      output ccl_mb_rip_h                      /* <bm1> */,
      output ccl_mb_rip_l                      /* <bm2> */,
      output ccl_mem_err_latch_l               /* <aa1> */,
      output ccl_mem_store_req_h               /* <ep1> */,
      output ccl_mem_store_req_l               /* <dl1> */,
      output ccl_mix_mb_sel_h                  /* <cf2> */,
      output ccl_odd_wc_par_h                  /* <dr2> */,
      output ccl_op_load_h                     /* <ec1> */,
      output ccl_op_load_l                     /* <cm1> */,
      output ccl_ram_req_l                     /* <bp2> */,
      output ccl_req_ctr_en_l                  /* <em2> */,
      output ccl_stSlres_intr_a_h              /* <cn1> */,
      output ccl_start_mem_l                   /* <de2> */,
      output ccl_wcEq0_in_h                    /* <cl1> */,
      output ccl_wcEq0_in_l                    /* <af2> */,
      output ccl_wcEq0_l                       /* <cl2> */,
      output ccl_wcEq1_h                       /* <fr2> */,
      output ccl_wcEq2_h                       /* <fr1> */,
      output ccl_wcEq3_h                       /* <fs1> */,
      output ccl_wc_ge4_l                      /* <ed1> */,
      output ccl_wd_taken_h                    /* <bu2> */,
      output ccl_zero_fill_h                   /* <ej2> */,
      output ccl_zero_fill_l                   /* <as1> */,
      input  ccw_act_flag_req_ena_h            /* <ca1> */,
      output ccw_buf_00_in_h                   /* <cm2> */,
      output ccw_buf_00_in_l                   /* <dr1> */,
      output ccw_buf_01_in_h                   /* <ds1> */,
      output ccw_buf_01_in_l                   /* <dp1> */,
      output ccw_buf_02_in_h                   /* <ea1> */,
      output ccw_buf_02_in_l                   /* <dm2> */,
      output ccw_buf_03_in_h                   /* <fs2> */,
      output ccw_buf_04_in_h                   /* <fp2> */,
      output ccw_buf_05_in_h                   /* <fn1> */,
      output ccw_buf_06_in_h                   /* <fm1> */,
      output ccw_buf_07_in_h                   /* <fj1> */,
      output ccw_buf_08_in_h                   /* <fk2> */,
      output ccw_buf_09_in_h                   /* <fk1> */,
      output ccw_buf_10_in_h                   /* <fl2> */,
      output ccw_buf_11_in_h                   /* <fl1> */,
      output ccw_buf_12_in_h                   /* <fm2> */,
      output ccw_buf_13_in_h                   /* <fp1> */,
      input  ccw_ccwf_req_ena_h                /* <cd2> */,
      input  ccw_cha_34_h                      /* <ep2> */,
      input  ccw_cha_35_h                      /* <en1> */,
      input  ccw_mem_adrEq0_l                  /* <bc1> */,
      input  ccw_mem_store_ena_h               /* <bv2> */,
      input  ccw_mix_00_h                      /* <cj2> */,
      input  ccw_mix_01_h                      /* <ck2> */,
      input  ccw_mix_02_h                      /* <ck1> */,
      input  ccw_mix_03_h                      /* <du2> */,
      input  ccw_mix_04_h                      /* <dn1> */,
      input  ccw_mix_05_h                      /* <dt2> */,
      input  ccw_mix_06_h                      /* <fd1> */,
      input  ccw_mix_07_h                      /* <fd2> */,
      input  ccw_mix_08_h                      /* <er1> */,
      input  ccw_mix_09_h                      /* <es2> */,
      input  ccw_mix_10_h                      /* <fe2> */,
      input  ccw_mix_11_h                      /* <ff2> */,
      input  ccw_mix_12_h                      /* <et2> */,
      input  ccw_mix_13_h                      /* <ev2> */,
      input  ccw_wd_ready_l                    /* <dj1> */,
      input  ch_ctom_l                         /* <cc1> */,
      input  ch_diag_04_l                      /* <da1> */,
      input  ch_diag_05_l                      /* <dc1> */,
      input  ch_diag_06_l                      /* <de1> */,
      input  ch_diag_read_a_l                  /* <dd2> */,
      input  ch_done_intr_h                    /* <an1> */,
      input  ch_done_intr_l                    /* <am2> */,
      input  ch_reset_intr_l                   /* <ch2> */,
      input  ch_reverse_h                      /* <cr1> */,
      input  ch_start_intr_l                   /* <cj1> */,
      input  ch_t0_l                           /* <as2> */,
      input  ch_t1_l                           /* <at2> */,
      input  ch_t2_l                           /* <au2> */,
      input  ch_t3_l                           /* <ap2> */,
      input  chan_adr_par_err_l                /* <ah2> */,
      input  chan_nxm_err_l                    /* <ak2> */,
      input  chan_par_err_l                    /* <bd2> */,
      input  clk_ccl_h                         /* <cr2> */,
      input  crc_act_ctr_0_h                   /* <em1> */,
      input  crc_act_ctr_1_h                   /* <dh2> */,
      input  crc_act_ctr_2_h                   /* <dj2> */,
      input  crc_act_ctr_2r_l                  /* <ef2> */,
      input  crc_mb_cyc_h                      /* <ce2> */,
      input  crc_mb_cyc_l                      /* <bl2> */,
      input  crc_ovn_err_in_h                  /* <eu2> */,
      input  crc_ram_adr_1r_h                  /* <br1> */,
      input  crc_ram_adr_2r_h                  /* <bn1> */,
      input  crc_ram_adr_4r_h                  /* <bp1> */,
      input  crc_ram_cyc_l                     /* <bf2> */,
      input  crc_req_d_h                       /* <dk1> */,
      input  crc_req_e_l                       /* <br2> */,
      input  crc_reset_l                       /* <ar2> */,
      input  crc_reverse_in_h                  /* <el2> */,
      input  crc_rh20_err_in_h                 /* <fe1> */,
      input  crc_short_wc_err_h                /* <es1> */,
      input  crc_wr_ram_l                      /* <ad2> */,
      input  csh_chan_cyc_a_h                  /* <cs1> */,
      output ebus_d00_e_h                      /* <dp2> */,
      output ebus_d02_e_h                      /* <ed2> */,
      output ebus_d03_e_h                      /* <cv2> */,
      input  mr_reset_05_h                     /* <al2> */
);

`include "ccl11nets.svh"

endmodule	// ccl11
