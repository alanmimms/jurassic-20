module cha;
`include "cha.svh"
endmodule	// cha
