module mtr;
`include "mtr.svh"
endmodule	// mtr
