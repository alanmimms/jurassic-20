module cac;
`include "cac.svh"
endmodule	// cac
