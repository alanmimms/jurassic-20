module mbz;
`include "mbz.svh"
endmodule	// mbz
