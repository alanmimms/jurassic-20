module mb015(
  /* <fc1> */ input  ar_06_a_h,
  /* <fd1> */ input  ar_07_a_h,
  /* <eu2> */ input  ar_08_a_h,
  /* <ev2> */ input  ar_09_a_h,
  /* <cv2> */ input  ar_10_a_h,
  /* <bu2> */ input  ar_11_a_h,
  /* <dd2> */ input  ar_24_a_h,
  /* <cs2> */ input  ar_25_a_h,
  /* <bp1> */ input  ar_26_a_h,
  /* <bj2> */ input  ar_27_a_h,
  /* <bm2> */ input  ar_28_a_h,
  /* <bf1> */ input  ar_29_a_h,
  /* <er2> */ input  cache_data_06_a_h,
  /* <ef1> */ input  cache_data_07_a_h,
  /* <ff2> */ input  cache_data_08_a_h,
  /* <er1> */ input  cache_data_09_a_h,
  /* <cr1> */ input  cache_data_10_a_h,
  /* <cm2> */ input  cache_data_11_a_h,
  /* <dk2> */ input  cache_data_24_a_h,
  /* <dk1> */ input  cache_data_25_a_h,
  /* <am1> */ input  cache_data_26_a_h,
  /* <ak1> */ input  cache_data_27_a_h,
  /* <ar1> */ input  cache_data_28_a_h,
  /* <ap1> */ input  cache_data_29_a_h,
  /* <cj1> */ input  cbus_d06_re_h,
  /* <ee1> */ output cbus_d06_te_h,
  /* <cj2> */ input  cbus_d07_re_h,
  /* <ee2> */ output cbus_d07_te_h,
  /* <bs2> */ input  cbus_d08_re_h,
  /* <el2> */ output cbus_d08_te_h,
  /* <bc1> */ input  cbus_d09_re_h,
  /* <em1> */ output cbus_d09_te_h,
  /* <br1> */ input  cbus_d10_re_h,
  /* <df1> */ output cbus_d10_te_h,
  /* <bd2> */ input  cbus_d11_re_h,
  /* <dl2> */ output cbus_d11_te_h,
  /* <ch2> */ input  cbus_d24_re_h,
  /* <dn1> */ output cbus_d24_te_h,
  /* <cf1> */ input  cbus_d25_re_h,
  /* <dm2> */ output cbus_d25_te_h,
  /* <be2> */ input  cbus_d26_re_h,
  /* <ah2> */ output cbus_d26_te_h,
  /* <bj1> */ input  cbus_d27_re_h,
  /* <af2> */ output cbus_d27_te_h,
  /* <be1> */ input  cbus_d28_re_h,
  /* <aj2> */ output cbus_d28_te_h,
  /* <bl1> */ input  cbus_d29_re_h,
  /* <ak2> */ output cbus_d29_te_h,
  /* <fk1> */ input  ccl_ccw_buf_wr_l,
  /* <ae2> */ input  ccl_ch_buf_en_l,
  /* <es1> */ input  ccl_mix_mb_sel_h,
  /* <fl1> */ input  ccw_buf_06_in_h,
  /* <fm2> */ input  ccw_buf_07_in_h,
  /* <fh2> */ input  ccw_buf_08_in_h,
  /* <fj2> */ input  ccw_buf_09_in_h,
  /* <cl2> */ input  ccw_buf_10_in_h,
  /* <cl1> */ input  ccw_buf_11_in_h,
  /* <ck2> */ input  ccw_buf_24_in_h,
  /* <ck1> */ input  ccw_buf_25_in_h,
  /* <at2> */ input  ccw_buf_26_in_h,
  /* <as1> */ input  ccw_buf_27_in_h,
  /* <ap2> */ input  ccw_buf_28_in_h,
  /* <am2> */ input  ccw_buf_29_in_h,
  /* <fk2> */ input  ccw_buf_adr_0_h,
  /* <fj1> */ input  ccw_buf_adr_1_h,
  /* <fl2> */ input  ccw_buf_adr_2_h,
  /* <fm1> */ input  ccw_buf_adr_3_h,
  /* <ek2> */ output ccw_mix_06_h,
  /* <eh2> */ output ccw_mix_07_h,
  /* <ff1> */ output ccw_mix_08_h,
  /* <es2> */ output ccw_mix_09_h,
  /* <cp2> */ output ccw_mix_10_h,
  /* <cn1> */ output ccw_mix_11_h,
  /* <dl1> */ output ccw_mix_24_h,
  /* <dh2> */ output ccw_mix_25_h,
  /* <al2> */ output ccw_mix_26_h,
  /* <al1> */ output ccw_mix_27_h,
  /* <as2> */ output ccw_mix_28_h,
  /* <ar2> */ output ccw_mix_29_h,
  /* <aj1> */ input  ch_buf_wr_04_l,
  /* <ep1> */ input  ch_buf_wr_1_l,
  /* <bd1> */ input  ch_reverse_h,
  /* <fs2> */ input  ch_t0_l,
  /* <af1> */ input  ch_t2_l,
  /* <cr2> */ input  clk_mb_06_h,
  /* <ek1> */ input  con_ki10_paging_mode_l,
  /* <dt2> */ input  crc_buf_mb_sel_h,
  /* <fu2> */ input  crc_cbus_out_hold_h,
  /* <fp2> */ input  crc_ch_buf_adr_0_h,
  /* <fr2> */ input  crc_ch_buf_adr_1_h,
  /* <fp1> */ input  crc_ch_buf_adr_2_h,
  /* <de1> */ input  crc_ch_buf_adr_3_h,
  /* <dj1> */ input  crc_ch_buf_adr_4_h,
  /* <de2> */ input  crc_ch_buf_adr_5_h,
  /* <ae1> */ input  crc_ch_buf_adr_6_h,
  /* <ad2> */ input  mb0_hold_in_h,
  /* <ad1> */ input  mb1_hold_in_h,
  /* <aa1> */ input  mb2_hold_in_h,
  /* <ac1> */ input  mb3_hold_in_h,
  /* <fc2> */ input  mb_06_h,
  /* <fd2> */ output mb_06_h,
  /* <ds2> */ output mb_06to11_par_odd_h,
  /* <dr2> */ output mb_07_h,
  /* <dp2> */ output mb_08_h,
  /* <dm1> */ output mb_09_h,
  /* <dr1> */ output mb_10_h,
  /* <dp1> */ output mb_11_h,
  /* <av2> */ output mb_24_h,
  /* <au2> */ output mb_24to29_par_odd_h,
  /* <ba1> */ output mb_25_h,
  /* <cd2> */ output mb_26_h,
  /* <cd1> */ output mb_27_h,
  /* <ca1> */ output mb_28_h,
  /* <bv2> */ output mb_29_h,
  /* <ej1> */ input  mb_in_sel_1_h,
  /* <el1> */ input  mb_in_sel_2_h,
  /* <ep2> */ input  mb_in_sel_4_h,
  /* <fr1> */ input  mb_sel_1_en_h,
  /* <ft2> */ input  mb_sel_2_en_h,
  /* <fv2> */ input  mb_sel_hold_h,
  /* <em2> */ input  mem_data_in_06_h,
  /* <ej2> */ input  mem_data_in_07_h,
  /* <ea1> */ input  mem_data_in_08_h,
  /* <dv2> */ input  mem_data_in_09_h,
  /* <cp1> */ input  mem_data_in_10_h,
  /* <cm1> */ input  mem_data_in_11_h,
  /* <dj2> */ input  mem_data_in_24_h,
  /* <df2> */ input  mem_data_in_25_h,
  /* <bm1> */ input  mem_data_in_26_h,
  /* <bk2> */ input  mem_data_in_27_h,
  /* <bl2> */ input  mem_data_in_28_h,
  /* <bk1> */ input  mem_data_in_29_h,
  /* <ed2> */ input  mem_to_c_en_l,
  /* <ed1> */ input  mem_to_c_sel_1_h,
  /* <ds1> */ input  mem_to_c_sel_2_h,
  /* <en1> */ output mem_to_cache_06_h,
  /* <ef2> */ output mem_to_cache_07_h,
  /* <ec1> */ output mem_to_cache_08_h,
  /* <du2> */ output mem_to_cache_09_h,
  /* <cf2> */ output mem_to_cache_10_h,
  /* <cc1> */ output mem_to_cache_11_h,
  /* <cs1> */ output mem_to_cache_24_h,
  /* <dd1> */ output mem_to_cache_25_h,
  /* <br2> */ output mem_to_cache_26_h,
  /* <bf2> */ output mem_to_cache_27_h,
  /* <bp2> */ output mem_to_cache_28_h,
  /* <bh2> */ output mem_to_cache_29_h,
  /* <fs1> */ input  nxm_any_l,
  /* <fe1> */ output pt_in_06_h,
  /* <fe2> */ output pt_in_07_h,
  /* <fa1> */ output pt_in_08_h,
  /* <et2> */ output pt_in_09_h,
  /* <dc1> */ output pt_in_10_h,
  /* <da1> */ output pt_in_11_h,
  /* <cu2> */ output pt_in_24_h,
  /* <ct2> */ output pt_in_25_h,
  /* <ce1> */ output pt_in_26_h,
  /* <ce2> */ output pt_in_27_h,
  /* <bs1> */ output pt_in_28_h,
  /* <bt2> */ output pt_in_29_h
);

`include "mb015nets.svh"

endmodule	// mb015
