module edp39(
  /* <cp2> */  input ad_28_h,
  /* <el2> */  input ad_29_h,
  /* <ck1> */ output ad_30_a_h,
  /* <cn1> */ output ad_30_a_l,
  /* <ep2> */ output ad_30_h,
  /* <at2> */ output ad_30to35Eq0_l,
  /* <dl1> */ output ad_31_h,
  /* <dr2> */ output ad_32_h,
  /* <dr1> */ output ad_33_h,
  /* <cf2> */ output ad_34_a_h,
  /* <cp1> */ output ad_34_h,
  /* <ce1> */ output ad_35_a_h,
  /* <el1> */ output ad_35_h,
  /* <am1> */ output ad_cg_30_h,
  /* <am2> */ output ad_cg_32_h,
  /* <aj1> */ output ad_cp_30_h,
  /* <af1> */ output ad_cp_32_h,
  /* <cu2> */ output ad_cry_31_h,
  /* <ct2> */ output ad_cry_31_l,
  /* <al1> */  input ad_cry_36_b_h,
  /* <cd1> */  input ad_cry_Ng02_a_h,
  /* <cv2> */ output ad_ex_28_h,
  /* <cr1> */ output ad_ex_29_h,
  /* <cl2> */ output ad_overflow_30_l,
  /* <ep1> */  input adx_00_h,
  /* <es2> */  input adx_29_h,
  /* <cf1> */ output adx_30_a_h,
  /* <cj2> */ output adx_30_h,
  /* <dk1> */ output adx_34_h,
  /* <es1> */ output adx_35_h,
  /* <al2> */ output adx_cg_30_h,
  /* <ak2> */ output adx_cg_33_h,
  /* <ae1> */ output adx_cp_30_h,
  /* <af2> */ output adx_cp_33_h,
  /* <fr2> */  input apr_fm_adr_10_h,
  /* <fp2> */  input apr_fm_adr_1_h,
  /* <fs1> */  input apr_fm_adr_2_h,
  /* <fn1> */  input apr_fm_adr_4_h,
  /* <fr1> */  input apr_fm_block_1_h,
  /* <fm1> */  input apr_fm_block_2_h,
  /* <fp1> */  input apr_fm_block_4_h,
  /* <fj2> */ output ar_30_a_h,
  /* <ft2> */ output ar_30_b_h,
  /* <fs2> */ output ar_30_c_h,
  /* <dm2> */ output ar_30_d_h,
  /* <bk2> */ output ar_30_h,
  /* <fc1> */ output ar_31_a_h,
  /* <fu2> */ output ar_31_b_h,
  /* <fv2> */ output ar_31_c_h,
  /* <bl2> */ output ar_31_h,
  /* <ff2> */ output ar_32_a_h,
  /* <cl1> */ output ar_32_b_h,
  /* <ch2> */ output ar_32_c_h,
  /* <eu2> */ output ar_33_a_h,
  /* <ck2> */ output ar_33_b_h,
  /* <cm1> */ output ar_33_c_h,
  /* <ev2> */ output ar_34_a_h,
  /* <fk1> */ output ar_34_b_h,
  /* <fk2> */ output ar_34_c_h,
  /* <et2> */ output ar_35_a_h,
  /* <fl2> */ output ar_35_b_h,
  /* <fl1> */ output ar_35_c_h,
  /* <em2> */  input armm_30_h,
  /* <ea1> */  input armm_31_h,
  /* <ee1> */  input armm_32_h,
  /* <dd2> */  input armm_33_h,
  /* <de1> */  input armm_34_h,
  /* <ef2> */  input armm_35_h,
  /* <bk1> */  input arx_00_h,
  /* <bl1> */  input arx_01_h,
  /* <as2> */ output arx_30_a_h,
  /* <br2> */ output arx_30_b_h,
  /* <ej2> */ output arx_30_h,
  /* <as1> */ output arx_31_a_h,
  /* <cm2> */ output arx_31_b_h,
  /* <bd2> */ output arx_31_h,
  /* <dc1> */ output arx_32_h,
  /* <aj2> */ output arx_33_h,
  /* <ac1> */ output arx_34_h,
  /* <aa1> */ output arx_35_h,
  /* <ej1> */  input arx_36_h,
  /* <bd1> */  input arx_37_h,
  /* <bm2> */ output br_30_a_h,
  /* <bm1> */  input brx_00_h,
  /* <be2> */ output brx_30_h,
  /* <be1> */  input brx_36_h,
  /* <em1> */  input cache_data_30_b_h,
  /* <ed2> */  input cache_data_31_b_h,
  /* <ee2> */  input cache_data_32_b_h,
  /* <dd1> */  input cache_data_33_b_h,
  /* <dl2> */  input cache_data_34_b_h,
  /* <cc1> */  input cache_data_35_b_h,
  /* <cr2> */  input clk_edp_30_h,
  /* <ce2> */  input con_fm_write_18to35_l,
  /* <ar1> */  input cram_Nr_30_h,
  /* <ap1> */  input cram_Nr_31_h,
  /* <ba1> */  input cram_Nr_32_h,
  /* <ap2> */  input cram_Nr_33_h,
  /* <av2> */  input cram_Nr_34_h,
  /* <au2> */  input cram_Nr_35_h,
  /* <an1> */  input cram_ad_boole_30_h,
  /* <ad2> */  input cram_ad_sel_1_30_h,
  /* <ah2> */  input cram_ad_sel_2_30_h,
  /* <ae2> */  input cram_ad_sel_4_30_h,
  /* <ad1> */  input cram_ad_sel_8_30_h,
  /* <bn1> */  input cram_ada_dis_30_h,
  /* <bj1> */  input cram_ada_sel_1_30_h,
  /* <bf2> */  input cram_ada_sel_2_30_h,
  /* <bt2> */  input cram_adb_sel_1_30_h,
  /* <bt1> */  input cram_adb_sel_1_30_h,
  /* <bs1> */  input cram_adb_sel_2_30_h,
  /* <er1> */  input cram_arm_sel_4_a_h,
  /* <ff1> */  input cram_arxm_sel_4_06_h,
  /* <dj2> */  input cram_br_load_a_h,
  /* <ar2> */  input cram_brx_load_a_h,
  /* <fe2> */  input ctl_ad_to_ebus_r_h,
  /* <ak1> */  input ctl_adx_cry_36_h,
  /* <eh2> */  input ctl_arr_clr_h,
  /* <ek2> */  input ctl_arr_load_a_l,
  /* <dh2> */  input ctl_arr_load_b_l,
  /* <en1> */  input ctl_arr_sel_1_h,
  /* <ek1> */  input ctl_arr_sel_2_h,
  /* <br1> */  input ctl_arx_load_h,
  /* <fj1> */  input ctl_arxr_sel_1_h,
  /* <fd2> */  input ctl_arxr_sel_2_h,
  /* <bu2> */  input ctl_mq_sel_1_h,
  /* <bv2> */  input ctl_mq_sel_2_h,
  /* <dn1> */  input ctl_mqm_en_h,
  /* <dj1> */  input ctl_mqm_sel_1_h,
  /* <dm1> */  input ctl_mqm_sel_2_h,
  /* <fd1> */  input diag_04_a_h,
  /* <fa1> */  input diag_05_a_h,
  /* <fe1> */  input diag_06_a_h,
  /* <ef1> */  input diag_read_func_12x_h,
  /* <dv2> */ output ebus_d30_e_h,
  /* <ds2> */ output ebus_d31_e_h,
  /* <dt2> */ output ebus_d32_e_h,
  /* <dp1> */ output ebus_d33_e_h,
  /* <dp2> */ output ebus_d34_e_h,
  /* <du2> */ output ebus_d35_e_h,
  /* <fm2> */ output edp_fm_parity_30to35_h,
  /* <cj1> */  input mq_00_h,
  /* <cs2> */  input mq_28_h,
  /* <cd2> */ output mq_30_h,
  /* <cs1> */ output mq_34_h,
  /* <df1> */ output mq_35_h,
  /* <ed1> */  input sh_30_h,
  /* <ec1> */  input sh_31_h,
  /* <ds1> */  input sh_32_h,
  /* <da1> */  input sh_33_h,
  /* <de2> */  input sh_34_h,
  /* <ca1> */  input sh_35_h,
  /* <bj2> */  input vma_held_or_pc_30_h,
  /* <bh2> */  input vma_held_or_pc_31_h,
  /* <bf1> */  input vma_held_or_pc_32_h,
  /* <bp2> */  input vma_held_or_pc_33_h,
  /* <bp1> */  input vma_held_or_pc_34_h,
  /* <bc1> */  input vma_held_or_pc_35_h
);

`include "edp39.svh"

endmodule	// edp39
