module edp49(
  /* <cp2> */ input  ad_10_h,
  /* <el2> */ input  ad_11_h,
  /* <ck1> */ output ad_12_a_h,
  /* <cn1> */ output ad_12_a_l,
  /* <ep2> */ output ad_12_h,
  /* <at2> */ output ad_12to17Eq0_l,
  /* <dl1> */ output ad_13_h,
  /* <dr2> */ output ad_14_h,
  /* <dr1> */ output ad_15_h,
  /* <cf2> */ output ad_16_a_h,
  /* <cp1> */ output ad_16_h,
  /* <ce1> */ output ad_17_a_h,
  /* <el1> */ output ad_17_h,
  /* <ep1> */ input  ad_18_h,
  /* <am1> */ output ad_cg_12_h,
  /* <am2> */ output ad_cg_14_h,
  /* <aj1> */ output ad_cp_12_h,
  /* <af1> */ output ad_cp_14_h,
  /* <cu2> */ output ad_cry_13_h,
  /* <ct2> */ output ad_cry_13_l,
  /* <al1> */ input  ad_cry_18_h,
  /* <cv2> */ output ad_ex_10_h,
  /* <cr1> */ output ad_ex_11_h,
  /* <cl2> */ output ad_overflow_12_l,
  /* <es2> */ input  adx_11_h,
  /* <cf1> */ output adx_12_a_h,
  /* <cj2> */ output adx_12_h,
  /* <dk1> */ output adx_16_h,
  /* <es1> */ output adx_17_h,
  /* <cj1> */ input  adx_18_h,
  /* <al2> */ output adx_cg_12_h,
  /* <ak2> */ output adx_cg_15_h,
  /* <ae1> */ output adx_cp_12_h,
  /* <af2> */ output adx_cp_15_h,
  /* <ak1> */ input  adx_cry_18_h,
  /* <fr2> */ input  apr_fm_adr_10_h,
  /* <fp2> */ input  apr_fm_adr_1_h,
  /* <fs1> */ input  apr_fm_adr_2_h,
  /* <fn1> */ input  apr_fm_adr_4_h,
  /* <fr1> */ input  apr_fm_block_1_h,
  /* <fm1> */ input  apr_fm_block_2_h,
  /* <fp1> */ input  apr_fm_block_4_h,
  /* <fj2> */ output ar_12_a_h,
  /* <ft2> */ output ar_12_b_h,
  /* <fs2> */ output ar_12_c_h,
  /* <dm2> */ output ar_12_d_h,
  /* <bk2> */ output ar_12_h,
  /* <fc1> */ output ar_13_a_h,
  /* <fu2> */ output ar_13_b_h,
  /* <fv2> */ output ar_13_c_h,
  /* <bl2> */ output ar_13_h,
  /* <ff2> */ output ar_14_a_h,
  /* <cl1> */ output ar_14_b_h,
  /* <ch2> */ output ar_14_c_h,
  /* <eu2> */ output ar_15_a_h,
  /* <ck2> */ output ar_15_b_h,
  /* <cm1> */ output ar_15_c_h,
  /* <ev2> */ output ar_16_a_h,
  /* <fk1> */ output ar_16_b_h,
  /* <fk2> */ output ar_16_c_h,
  /* <et2> */ output ar_17_a_h,
  /* <fl2> */ output ar_17_b_h,
  /* <fl1> */ output ar_17_c_h,
  /* <bk1> */ input  ar_18_h,
  /* <bl1> */ input  ar_19_h,
  /* <em2> */ input  armm_12_h,
  /* <ea1> */ input  armm_13_h,
  /* <ee1> */ input  armm_14_h,
  /* <dd2> */ input  armm_15_h,
  /* <de1> */ input  armm_16_h,
  /* <ef2> */ input  armm_17_h,
  /* <as2> */ output arx_12_a_h,
  /* <br2> */ output arx_12_b_h,
  /* <ej2> */ output arx_12_h,
  /* <as1> */ output arx_13_a_h,
  /* <cm2> */ output arx_13_b_h,
  /* <bd2> */ output arx_13_h,
  /* <dc1> */ output arx_14_h,
  /* <aj2> */ output arx_15_h,
  /* <ac1> */ output arx_16_h,
  /* <aa1> */ output arx_17_h,
  /* <ej1> */ input  arx_18_h,
  /* <bd1> */ input  arx_19_h,
  /* <bm2> */ output br_12_a_h,
  /* <bm1> */ input  br_18_a_h,
  /* <be2> */ output brx_12_h,
  /* <be1> */ input  brx_18_h,
  /* <em1> */ input  cache_data_12_b_h,
  /* <ed2> */ input  cache_data_13_b_h,
  /* <ee2> */ input  cache_data_14_b_h,
  /* <dd1> */ input  cache_data_15_b_h,
  /* <dl2> */ input  cache_data_16_b_h,
  /* <cc1> */ input  cache_data_17_b_h,
  /* <cr2> */ input  clk_edp_12_h,
  /* <ce2> */ input  con_fm_write_00to17_l,
  /* <ar1> */ input  cram_Nr_12_h,
  /* <ap1> */ input  cram_Nr_13_h,
  /* <ba1> */ input  cram_Nr_14_h,
  /* <ap2> */ input  cram_Nr_15_h,
  /* <av2> */ input  cram_Nr_16_h,
  /* <au2> */ input  cram_Nr_17_h,
  /* <an1> */ input  cram_ad_boole_12_h,
  /* <ad2> */ input  cram_ad_sel_1_12_h,
  /* <ah2> */ input  cram_ad_sel_2_12_h,
  /* <ae2> */ input  cram_ad_sel_4_12_h,
  /* <ad1> */ input  cram_ad_sel_8_12_h,
  /* <bn1> */ input  cram_ada_dis_12_h,
  /* <bj1> */ input  cram_ada_sel_1_12_h,
  /* <bf2> */ input  cram_ada_sel_2_12_h,
  /* <bt2> */ input  cram_adb_sel_1_12_h,
  /* <bt1> */ input  cram_adb_sel_1_12_h,
  /* <bs1> */ input  cram_adb_sel_2_12_h,
  /* <ff1> */ input  cram_arxm_sel_4_00_h,
  /* <dj2> */ input  cram_br_load_a_h,
  /* <ar2> */ input  cram_brx_load_a_h,
  /* <fe2> */ input  ctl_ad_to_ebus_l_h,
  /* <ek2> */ input  ctl_ar_09to17_load_l,
  /* <dh2> */ input  ctl_ar_09to17_load_l,
  /* <eh2> */ input  ctl_ar_12to17_clr_h,
  /* <en1> */ input  ctl_arl_sel_1_h,
  /* <ek1> */ input  ctl_arl_sel_2_h,
  /* <er1> */ input  ctl_arl_sel_4_h,
  /* <br1> */ input  ctl_arx_load_h,
  /* <fj1> */ input  ctl_arxl_sel_1_h,
  /* <fd2> */ input  ctl_arxl_sel_2_h,
  /* <bu2> */ input  ctl_mq_sel_1_h,
  /* <bv2> */ input  ctl_mq_sel_2_h,
  /* <dn1> */ input  ctl_mqm_en_h,
  /* <dj1> */ input  ctl_mqm_sel_1_h,
  /* <dm1> */ input  ctl_mqm_sel_2_h,
  /* <fd1> */ input  diag_04_a_h,
  /* <fa1> */ input  diag_05_a_h,
  /* <fe1> */ input  diag_06_a_h,
  /* <ef1> */ input  diag_read_func_12x_h,
  /* <dv2> */ output ebus_d12_e_h,
  /* <ds2> */ output ebus_d13_e_h,
  /* <dt2> */ output ebus_d14_e_h,
  /* <dp1> */ output ebus_d15_e_h,
  /* <dp2> */ output ebus_d16_e_h,
  /* <du2> */ output ebus_d17_e_h,
  /* <fm2> */ output edp_fm_parity_12to17_h,
  /* <cs2> */ input  mq_10_h,
  /* <cd2> */ output mq_12_h,
  /* <cs1> */ output mq_16_h,
  /* <df1> */ output mq_17_h,
  /* <cd1> */ input  mq_18_h,
  /* <ed1> */ input  sh_12_h,
  /* <ec1> */ input  sh_13_h,
  /* <ds1> */ input  sh_14_h,
  /* <da1> */ input  sh_15_h,
  /* <de2> */ input  sh_16_h,
  /* <ca1> */ input  sh_17_h,
  /* <bj2> */ input  vma_held_or_pc_12_h,
  /* <bh2> */ input  vma_held_or_pc_13_h,
  /* <bf1> */ input  vma_held_or_pc_14_h,
  /* <bp2> */ input  vma_held_or_pc_15_h,
  /* <bp1> */ input  vma_held_or_pc_16_h,
  /* <bc1> */ input  vma_held_or_pc_17_h
);

`include "edp49nets.svh"

endmodule	// edp49
