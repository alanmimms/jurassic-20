module tapped_delay_20_2(input bit in, output bit t1,t2,t3,t4,t5,t6,t7,t8,t9, out);
  assign t1 = in;
  assign t2 = in;
  assign t3 = in;
  assign t4 = in;
  assign t5 = in;
  assign t6 = in;
  assign t7 = in;
  assign t8 = in;
  assign t9 = in;
  assign out = in;
endmodule // tapped_delay_20_2
