module edp;
`include "edp.svh"
endmodule	// edp
