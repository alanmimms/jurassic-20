module ccl;
`include "ccl.svh"
endmodule	// ccl
