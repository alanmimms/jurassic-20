module scd54(
  /* <bd2> */  input ad_cry_01_l,
  /* <ar2> */  input ad_cry_Ng02_a_l,
  /* <bd1> */  input ad_overflow_00_l,
  /* <dm1> */  input ar_00_d_h,
  /* <fu2> */  input ar_01_c_h,
  /* <fr2> */  input ar_02_c_h,
  /* <ff1> */  input ar_03_c_h,
  /* <fk2> */  input ar_04_c_h,
  /* <dh2> */  input ar_05_c_h,
  /* <dl1> */  input ar_06_c_h,
  /* <ev2> */  input ar_07_c_h,
  /* <de2> */  input ar_08_c_h,
  /* <df2> */  input ar_09_c_h,
  /* <ds1> */  input ar_10_c_h,
  /* <dm2> */  input ar_11_c_h,
  /* <fd2> */  input ar_18_c_h,
  /* <fc1> */  input ar_28_c_h,
  /* <ff2> */  input ar_29_c_h,
  /* <fd1> */  input ar_30_c_h,
  /* <fj2> */  input ar_31_c_h,
  /* <ee1> */  input ar_32_c_h,
  /* <cv2> */  input ar_33_c_h,
  /* <ef1> */  input ar_34_c_h,
  /* <cs1> */  input ar_35_c_h,
  /* <dj1> */ output armm_00_h,
  /* <dd1> */ output armm_01_h,
  /* <dl2> */ output armm_02_h,
  /* <df1> */ output armm_03_h,
  /* <dk1> */ output armm_04_h,
  /* <dc1> */ output armm_05_h,
  /* <cm1> */ output armm_06_h,
  /* <cl2> */ output armm_07_h,
  /* <ck1> */ output armm_08_h,
  /* <cr2> */  input clk3_scd_h,
  /* <af2> */  input clk_mb_xfer_l,
  /* <ba1> */  input con_clr_private_instr_h,
  /* <ac1> */  input con_condSlad_flags_h,
  /* <es2> */  input con_condSlfe_shrt_h,
  /* <br1> */  input con_condSlpcfGETSNr_h,
  /* <cs2> */  input con_cond_en_30to37_l,
  /* <er2> */  input con_cond_instr_abort_h,
  /* <bf1> */  input con_fm_xfer_l,
  /* <ad2> */  input con_nicond_trap_en_h,
  /* <ch2> */  input con_pcPl1_inh_l,
  /* <bu2> */  input con_pi_cycle_a_l,
  /* <bf2> */  input con_trap_en_a_h,
  /* <es1> */  input cram_Nr_00_h,
  /* <ft2> */  input cram_Nr_01_h,
  /* <fp2> */  input cram_Nr_02_h,
  /* <fe1> */  input cram_Nr_03_h,
  /* <fl2> */  input cram_Nr_04_h,
  /* <dd2> */  input cram_Nr_05_h,
  /* <cu2> */  input cram_Nr_06_h,
  /* <dr1> */  input cram_Nr_07_h,
  /* <cp1> */  input cram_Nr_08_h,
  /* <cp2> */  input cram_cond_03_a_h,
  /* <ed1> */  input cram_cond_04_a_h,
  /* <ct2> */  input cram_cond_05_a_h,
  /* <eu2> */  input cram_scad_1_h,
  /* <dr2> */  input cram_scad_2_h,
  /* <dp1> */  input cram_scad_4_h,
  /* <fk1> */  input cram_scada_en_l,
  /* <fl1> */  input cram_scada_sel_1_h,
  /* <fj1> */  input cram_scada_sel_2_h,
  /* <fs2> */  input cram_scadb_sel_1_h,
  /* <fm2> */  input cram_scadb_sel_2_h,
  /* <fa1> */  input cram_scm_sel_2_h,
  /* <de1> */  input cram_shNgarmm_sel_1_h,
  /* <da1> */  input cram_shNgarmm_sel_2_h,
  /* <cj2> */  input cram_vma_sel_2_a_h,
  /* <br2> */  input ctl1_condSlarGETSexp_h,
  /* <aa1> */  input ctl1_specSlclr_fpd_h,
  /* <bj2> */  input ctl1_specSlflag_ctl_h,
  /* <fe2> */  input ctl1_specSlscm_alt_h,
  /* <et2> */  input ctl_dispSlnicond_h,
  /* <ae2> */  input ctl_specSlsave_flags_l,
  /* <cf2> */  input diag_04_a_h,
  /* <ce2> */  input diag_05_a_h,
  /* <bp1> */  input diag_06_a_h,
  /* <bn1> */  input diag_read_func_13x_l,
  /* <ce1> */ output ebus_d02_e_h,
  /* <cf1> */ output ebus_d03_e_h,
  /* <cd1> */ output ebus_d04_e_h,
  /* <cc1> */ output ebus_d05_e_h,
  /* <ca1> */ output ebus_d06_e_h,
  /* <ea1> */ output ebus_d07_e_h,
  /* <dt2> */ output ebus_d08_e_h,
  /* <dv2> */ output ebus_d09_e_h,
  /* <ds2> */ output ebus_d10_e_h,
  /* <du2> */ output ebus_d11_e_h,
  /* <bl2> */  input mcl6_paged_fetch_l,
  /* <bl1> */  input mr_reset_01_h,
  /* <ck2> */  input pi2_pi1_a_l,
  /* <cm2> */  input pi2_pi2_a_l,
  /* <cl1> */  input pi2_pi4_a_l,
  /* <bp2> */  input pt_public_h,
  /* <bt2> */ output scd1_scadEq0_l,
  /* <fv2> */ output scd1_scad_sign_h,
  /* <ek1> */ output scd2_fe_sign_h,
  /* <ee2> */ output scd2_sc_04_h,
  /* <er1> */ output scd2_sc_05_h,
  /* <dj2> */ output scd2_sc_06_h,
  /* <dk2> */ output scd2_sc_07_h,
  /* <ed2> */ output scd2_sc_08_h,
  /* <ef2> */ output scd2_sc_09_h,
  /* <em2> */ output scd2_sc_36_to_63_h,
  /* <el2> */ output scd2_sc_DtgeDt_36_h,
  /* <ej1> */ output scd2_sc_sign_h,
  /* <bm2> */ output scd3_trap_mix_32_h,
  /* <cj1> */ output scd3_trap_mix_33_h,
  /* <bm1> */ output scd3_trap_mix_34_h,
  /* <cd2> */ output scd3_trap_mix_35_h,
  /* <bk2> */ output scd4_cry0_h,
  /* <bs1> */ output scd4_cry1_h,
  /* <as2> */ output scd4_div_chk_h,
  /* <bk1> */ output scd4_fov_h,
  /* <ap2> */ output scd4_fpd_h,
  /* <bs2> */ output scd4_fxu_h,
  /* <am2> */ output scd4_nicond_10_h,
  /* <ak2> */ output scd4_pcp_h,
  /* <bc1> */ output scd4_trap_req_1_h,
  /* <ad1> */ output scd4_trap_req_2_h,
  /* <bj1> */ output scd5_adr_brk_inh_h,
  /* <au2> */ output scd5_adr_brk_prevent_h,
  /* <aj2> */ output scd5_adr_brk_prevent_l,
  /* <av2> */ output scd5_kernelSluser_iot_h,
  /* <ah2> */ output scd5_private_instr_l,
  /* <dp2> */ output scd5_public_a_h,
  /* <cr1> */ output scd5_user_a_h,
  /* <be2> */ output scd5_user_iot_a_h,
  /* <bv2> */ output scd_kernel_mode_h,
  /* <ae1> */ output scd_public_a_l,
  /* <at2> */ output scd_user_a_l,
  /* <af1> */ output scd_user_iot_a_l,
  /* <al2> */ output vma_held_or_pc_00_h
);

`include "scd54nets.svh"

endmodule	// scd54
