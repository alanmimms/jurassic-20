module cac17(
  /* <cv2> */  input cache_adr_27_h,
  /* <da1> */  input cache_adr_28_h,
  /* <dp1> */  input cache_adr_29_h,
  /* <dv2> */  input cache_adr_30_h,
  /* <es1> */  input cache_adr_31_h,
  /* <cf1> */  input cache_adr_32_h,
  /* <ca1> */  input cache_adr_33_h,
  /* <bf1> */  input cache_adr_34_h,
  /* <br1> */  input cache_adr_35_h,
  /* <bs1> */  input cache_adr_35_l,
  /* <ff1> */ output cache_data_27_a_h,
  /* <fe2> */ output cache_data_27_b_h,
  /* <fe1> */ output cache_data_27_c_h,
  /* <ep2> */ output cache_data_28_a_h,
  /* <ep1> */ output cache_data_28_b_h,
  /* <er1> */ output cache_data_28_c_h,
  /* <es2> */ output cache_data_29_a_h,
  /* <eu2> */ output cache_data_29_b_h,
  /* <ev2> */ output cache_data_29_c_h,
  /* <df1> */ output cache_data_30_a_h,
  /* <df2> */ output cache_data_30_b_h,
  /* <de1> */ output cache_data_30_c_h,
  /* <dm1> */ output cache_data_31_a_h,
  /* <dm2> */ output cache_data_31_b_h,
  /* <dl2> */ output cache_data_31_c_h,
  /* <be2> */ output cache_data_32_a_h,
  /* <be1> */ output cache_data_32_b_h,
  /* <bf2> */ output cache_data_32_c_h,
  /* <bk1> */ output cache_data_33_a_h,
  /* <bl2> */ output cache_data_33_b_h,
  /* <bk2> */ output cache_data_33_c_h,
  /* <ar1> */ output cache_data_34_a_h,
  /* <ap2> */ output cache_data_34_b_h,
  /* <ar2> */ output cache_data_34_c_h,
  /* <bd2> */ output cache_data_35_a_h,
  /* <ba1> */ output cache_data_35_b_h,
  /* <bd1> */ output cache_data_35_c_h,
  /* <el1> */  input cache_wr_27_a_l,
  /* <ej1> */  input csh_0_00to17_sel_a_l,
  /* <ee1> */  input csh_1_00to17_sel_a_l,
  /* <bj2> */  input csh_2_00to17_sel_a_l,
  /* <bj1> */  input csh_3_00to17_sel_a_l,
  /* <dd1> */ output csh_par_bit_03_a_h,
  /* <fa1> */ output csh_par_bit_03_b_h,
  /* <fd1> */  input csh_par_bit_in_h,
  /* <fd2> */  input mem_to_cache_27_h,
  /* <er2> */  input mem_to_cache_28_h,
  /* <ff2> */  input mem_to_cache_29_h,
  /* <cm1> */  input mem_to_cache_30_h,
  /* <cp1> */  input mem_to_cache_31_h,
  /* <cl1> */  input mem_to_cache_32_h,
  /* <au2> */  input mem_to_cache_33_h,
  /* <av2> */  input mem_to_cache_34_h,
  /* <as2> */  input mem_to_cache_35_h
);

`include "cac17nets.svh"

endmodule	// cac17
