module edp41(
      output ad_22_h                           /* <cv2> */,
      output ad_23_h                           /* <cr1> */,
      output ad_24_a_h                         /* <ck1> */,
      output ad_24_a_l                         /* <cn1> */,
      output ad_24_h                           /* <ep2> */,
      output ad_24to29Eq0_l                    /* <at2> */,
      output ad_25_h                           /* <dl1> */,
      output ad_26_h                           /* <dr2> */,
      output ad_27_h                           /* <dr1> */,
      output ad_28_a_h                         /* <cf2> */,
      output ad_28_h                           /* <cp1> */,
      output ad_29_a_h                         /* <ce1> */,
      output ad_29_h                           /* <el1> */,
      input  ad_30_h                           /* <ep1> */,
      output ad_cg_24_h                        /* <am1> */,
      output ad_cg_26_h                        /* <am2> */,
      output ad_cp_24_h                        /* <aj1> */,
      output ad_cp_26_h                        /* <af1> */,
      output ad_cry_25_h                       /* <cu2> */,
      output ad_cry_25_l                       /* <ct2> */,
      input  ad_cry_30_h                       /* <al1> */,
      output ad_overflow_24_l                  /* <cl2> */,
      input  adx_23_h                          /* <es2> */,
      output adx_24_a_h                        /* <cf1> */,
      output adx_24_h                          /* <cj2> */,
      output adx_28_h                          /* <dk1> */,
      output adx_29_h                          /* <es1> */,
      input  adx_30_h                          /* <cj1> */,
      output adx_cg_24_h                       /* <al2> */,
      output adx_cg_27_h                       /* <ak2> */,
      output adx_cp_24_h                       /* <ae1> */,
      output adx_cp_27_h                       /* <af2> */,
      input  adx_cry_30_h                      /* <ak1> */,
      input  apr_fm_adr_10_h                   /* <fr2> */,
      input  apr_fm_adr_1_h                    /* <fp2> */,
      input  apr_fm_adr_2_h                    /* <fs1> */,
      input  apr_fm_adr_4_h                    /* <fn1> */,
      input  apr_fm_block_1_h                  /* <fr1> */,
      input  apr_fm_block_2_h                  /* <fm1> */,
      input  apr_fm_block_4_h                  /* <fp1> */,
      output ar_24_a_h                         /* <fj2> */,
      output ar_24_b_h                         /* <ft2> */,
      output ar_24_c_h                         /* <fs2> */,
      output ar_24_d_h                         /* <dm2> */,
      output ar_24_h                           /* <bk2> */,
      output ar_25_a_h                         /* <fc1> */,
      output ar_25_b_h                         /* <fu2> */,
      output ar_25_c_h                         /* <fv2> */,
      output ar_25_h                           /* <bl2> */,
      output ar_26_a_h                         /* <ff2> */,
      output ar_26_b_h                         /* <cl1> */,
      output ar_26_c_h                         /* <ch2> */,
      output ar_27_a_h                         /* <eu2> */,
      output ar_27_b_h                         /* <ck2> */,
      output ar_27_c_h                         /* <cm1> */,
      output ar_28_a_h                         /* <ev2> */,
      output ar_28_b_h                         /* <fk1> */,
      output ar_28_c_h                         /* <fk2> */,
      output ar_29_a_h                         /* <et2> */,
      output ar_29_b_h                         /* <fl2> */,
      output ar_29_c_h                         /* <fl1> */,
      input  ar_30_h                           /* <bk1> */,
      input  ar_31_h                           /* <bl1> */,
      input  armm_24_h                         /* <em2> */,
      input  armm_25_h                         /* <ea1> */,
      input  armm_26_h                         /* <ee1> */,
      input  armm_27_h                         /* <dd2> */,
      input  armm_28_h                         /* <de1> */,
      input  armm_29_h                         /* <ef2> */,
      output arx_24_a_h                        /* <as2> */,
      output arx_24_b_h                        /* <br2> */,
      output arx_24_h                          /* <ej2> */,
      output arx_25_a_h                        /* <as1> */,
      output arx_25_b_h                        /* <cm2> */,
      output arx_25_h                          /* <bd2> */,
      output arx_26_h                          /* <dc1> */,
      output arx_27_h                          /* <aj2> */,
      output arx_28_h                          /* <ac1> */,
      output arx_29_h                          /* <aa1> */,
      input  arx_30_h                          /* <ej1> */,
      input  arx_31_h                          /* <bd1> */,
      output br_24_a_h                         /* <bm2> */,
      input  br_30_a_h                         /* <bm1> */,
      output brx_24_h                          /* <be2> */,
      input  brx_30_h                          /* <be1> */,
      input  cache_data_24_b_h                 /* <em1> */,
      input  cache_data_25_b_h                 /* <ed2> */,
      input  cache_data_26_b_h                 /* <ee2> */,
      input  cache_data_27_b_h                 /* <dd1> */,
      input  cache_data_28_b_h                 /* <dl2> */,
      input  cache_data_29_b_h                 /* <cc1> */,
      input  clk_edp_24_h                      /* <cr2> */,
      input  con_fm_write_18to35_l             /* <ce2> */,
      input  cram_Nr_24_h                      /* <ar1> */,
      input  cram_Nr_25_h                      /* <ap1> */,
      input  cram_Nr_26_h                      /* <ba1> */,
      input  cram_Nr_27_h                      /* <ap2> */,
      input  cram_Nr_28_h                      /* <av2> */,
      input  cram_Nr_29_h                      /* <au2> */,
      input  cram_ad_boole_24_h                /* <an1> */,
      input  cram_ad_sel_1_24_h                /* <ad2> */,
      input  cram_ad_sel_2_24_h                /* <ah2> */,
      input  cram_ad_sel_4_24_h                /* <ae2> */,
      input  cram_ad_sel_8_24_h                /* <ad1> */,
      input  cram_ada_dis_24_h                 /* <bn1> */,
      input  cram_ada_sel_1_24_h               /* <bj1> */,
      input  cram_ada_sel_2_24_h               /* <bf2> */,
      input  cram_adb_sel_1_24_h               /* <bt2> */,
      input  cram_adb_sel_2_24_h               /* <bs1> */,
      input  cram_arm_sel_4_a_h                /* <er1> */,
      input  cram_arxm_sel_4_06_h              /* <ff1> */,
      input  cram_br_load_a_h                  /* <dj2> */,
      input  cram_brx_load_a_h                 /* <ar2> */,
      input  ctl_ad_to_ebus_r_h                /* <fe2> */,
      input  ctl_arr_clr_h                     /* <eh2> */,
      input  ctl_arr_load_a_l                  /* <ek2> */,
      input  ctl_arr_load_b_l                  /* <dh2> */,
      input  ctl_arr_sel_1_h                   /* <en1> */,
      input  ctl_arr_sel_2_h                   /* <ek1> */,
      input  ctl_arx_load_h                    /* <br1> */,
      input  ctl_arxr_sel_1_h                  /* <fj1> */,
      input  ctl_arxr_sel_2_h                  /* <fd2> */,
      input  ctl_mq_sel_1_h                    /* <bu2> */,
      input  ctl_mq_sel_2_h                    /* <bv2> */,
      input  ctl_mqm_en_h                      /* <dn1> */,
      input  ctl_mqm_sel_1_h                   /* <dj1> */,
      input  ctl_mqm_sel_2_h                   /* <dm1> */,
      input  diag_04_a_h                       /* <fd1> */,
      input  diag_05_a_h                       /* <fa1> */,
      input  diag_06_a_h                       /* <fe1> */,
      input  diag_read_func_12x_h              /* <ef1> */,
      output ebus_d24_e_h                      /* <dv2> */,
      output ebus_d25_e_h                      /* <ds2> */,
      output ebus_d26_e_h                      /* <dt2> */,
      output ebus_d27_e_h                      /* <dp1> */,
      output ebus_d28_e_h                      /* <dp2> */,
      output ebus_d29_e_h                      /* <du2> */,
      output edp_fm_parity_24to29_h            /* <fm2> */,
      input  mq_22_h                           /* <cs2> */,
      output mq_24_h                           /* <cd2> */,
      output mq_28_h                           /* <cs1> */,
      output mq_29_h                           /* <df1> */,
      input  mq_30_h                           /* <cd1> */,
      input  sh_24_h                           /* <ed1> */,
      input  sh_25_h                           /* <ec1> */,
      input  sh_26_h                           /* <ds1> */,
      input  sh_27_h                           /* <da1> */,
      input  sh_28_h                           /* <de2> */,
      input  sh_29_h                           /* <ca1> */,
      input  vma_held_or_pc_24_h               /* <bj2> */,
      input  vma_held_or_pc_25_h               /* <bh2> */,
      input  vma_held_or_pc_26_h               /* <bf1> */,
      input  vma_held_or_pc_27_h               /* <bp2> */,
      input  vma_held_or_pc_28_h               /* <bp1> */,
      input  vma_held_or_pc_29_h               /* <bc1> */
);

`include "edp41nets.svh"

endmodule	// edp41
