module cac19(
      input  cache_adr_27_h                    /* <cv2> */,
      input  cache_adr_28_h                    /* <da1> */,
      input  cache_adr_29_h                    /* <dp1> */,
      input  cache_adr_30_h                    /* <dv2> */,
      input  cache_adr_31_h                    /* <es1> */,
      input  cache_adr_32_h                    /* <cf1> */,
      input  cache_adr_33_h                    /* <ca1> */,
      input  cache_adr_34_h                    /* <bf1> */,
      input  cache_adr_35_h                    /* <br1> */,
      input  cache_adr_35_l                    /* <bs1> */,
      output cache_data_18_a_h                 /* <ff1> */,
      output cache_data_18_b_h                 /* <fe2> */,
      output cache_data_18_c_h                 /* <fe1> */,
      output cache_data_19_a_h                 /* <ep2> */,
      output cache_data_19_b_h                 /* <ep1> */,
      output cache_data_19_c_h                 /* <er1> */,
      output cache_data_20_a_h                 /* <es2> */,
      output cache_data_20_b_h                 /* <eu2> */,
      output cache_data_20_c_h                 /* <ev2> */,
      output cache_data_21_a_h                 /* <df1> */,
      output cache_data_21_b_h                 /* <df2> */,
      output cache_data_21_c_h                 /* <de1> */,
      output cache_data_22_a_h                 /* <dm1> */,
      output cache_data_22_b_h                 /* <dm2> */,
      output cache_data_22_c_h                 /* <dl2> */,
      output cache_data_23_a_h                 /* <be2> */,
      output cache_data_23_b_h                 /* <be1> */,
      output cache_data_23_c_h                 /* <bf2> */,
      output cache_data_24_a_h                 /* <bk1> */,
      output cache_data_24_b_h                 /* <bl2> */,
      output cache_data_24_c_h                 /* <bk2> */,
      output cache_data_25_a_h                 /* <ar1> */,
      output cache_data_25_b_h                 /* <ap2> */,
      output cache_data_25_c_h                 /* <ar2> */,
      output cache_data_26_a_h                 /* <bd2> */,
      output cache_data_26_b_h                 /* <ba1> */,
      output cache_data_26_c_h                 /* <bd1> */,
      input  cache_wr_18_a_l                   /* <el1> */,
      input  csh_0_00to17_sel_a_l              /* <ej1> */,
      input  csh_1_00to17_sel_a_l              /* <ee1> */,
      input  csh_2_00to17_sel_a_l              /* <bj2> */,
      input  csh_2_0to17_sel_a_l               /* <as1> */,
      input  csh_3_00to17_sel_a_l              /* <bj1> */,
      input  csh_en_csh_data_l                 /* <ck1> */,
      output csh_par_bit_02_a_h                /* <dd1> */,
      output csh_par_bit_02_b_h                /* <fa1> */,
      input  csh_par_bit_in_h                  /* <fd1> */,
      input  mem_to_cache_18_h                 /* <fd2> */,
      input  mem_to_cache_19_h                 /* <er2> */,
      input  mem_to_cache_20_h                 /* <ff2> */,
      input  mem_to_cache_21_h                 /* <cm1> */,
      input  mem_to_cache_22_h                 /* <cp1> */,
      input  mem_to_cache_23_h                 /* <cl1> */,
      input  mem_to_cache_24_h                 /* <au2> */,
      input  mem_to_cache_25_h                 /* <av2> */,
      input  mem_to_cache_26_h                 /* <as2> */
);

`include "cac19nets.svh"

endmodule	// cac19
