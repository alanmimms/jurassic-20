module mb0;
`include "mb0.svh"
endmodule	// mb0
