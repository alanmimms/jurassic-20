module csh23(
      input  a_change_coming_in_l              /* <bc1> */,
      input  apr6_ebox_cca_l                   /* <da1> */,
      input  apr6_ebox_era_l                   /* <ba1> */,
      input  apr6_ebox_load_reg_l              /* <ds1> */,
      input  apr6_ebox_read_reg_h              /* <aj1> */,
      input  apr6_ebox_read_reg_l              /* <av2> */,
      input  apr6_ebox_sbus_diag_h             /* <ak1> */,
      input  apr_ebox_sbus_diag_l              /* <dk1> */,
      input  apr_en_refill_ram_wr_h            /* <fr1> */,
      input  cache_to_mb_t4_l                  /* <ef2> */,
      input  ccl_chan_req_h                    /* <fe1> */,
      input  ccl_chan_req_l                    /* <fl1> */,
      input  ccl_chan_to_mem_h                 /* <af1> */,
      input  ccl_chan_to_mem_l                 /* <dt2> */,
      input  chan_read_h                       /* <ce1> */,
      input  clk1_csh_h                        /* <cr2> */,
      input  clk3_ebox_sync_d_l                /* <ej2> */,
      input  clk4_ebox_cyc_abort_h             /* <fa1> */,
      input  clk4_ebox_req_h                   /* <fh2> */,
      input  clk4_ebox_req_l                   /* <ee1> */,
      input  con_ki10_paging_mode_h            /* <at2> */,
      input  core_busy_h                       /* <ec1> */,
      input  core_busy_l                       /* <fv2> */,
      output csh1_cca_cyc_l                    /* <ap2> */,
      output csh1_cca_req_grant_h              /* <eu2> */,
      output csh1_chan_req_grant_h             /* <ev2> */,
      output csh1_ebox_cca_grant_h             /* <ca1> */,
      output csh1_ebox_era_grant_h             /* <aa1> */,
      output csh1_ebox_req_grant_a_l           /* <es1> */,
      output csh1_ebox_req_grant_h             /* <ek2> */,
      output csh1_mb_cyc_l                     /* <bp2> */,
      output csh1_mb_req_grant_l               /* <et2> */,
      output csh1_pgrf_cyc_a_h                 /* <bk2> */,
      output csh1_pgrf_cyc_a_l                 /* <bj2> */,
      output csh1_ready_to_go_h                /* <fm1> */,
      output csh1_ready_to_go_l                /* <cc1> */,
      output csh2_e_cache_wr_cyc_h             /* <em2> */,
      output csh2_e_core_rd_rq_b_l             /* <ea1> */,
      output csh2_e_core_rd_rq_l               /* <fs2> */,
      output csh2_ebox_retry_req_l             /* <as1> */,
      output csh2_mbox_resp_in_h               /* <bd1> */,
      output csh2_one_word_rd_h                /* <bk1> */,
      output csh2_one_word_rd_l                /* <be2> */,
      output csh2_rd_pause_2nd_half_l          /* <dp2> */,
      output csh3_adr_pma_en_h                 /* <ep2> */,
      output csh3_adr_ready_l                  /* <fj1> */,
      output csh3_any_val_hold_a_h             /* <fr2> */,
      output csh3_any_val_hold_in_h            /* <ff1> */,
      output csh3_gate_vma_27to33_h            /* <ep1> */,
      output csh3_match_hold_1_in_h            /* <br2> */,
      output csh3_match_hold_2_in_h            /* <bu2> */,
      output csh3_mb_wr_rq_clr_nxt_l           /* <fm2> */,
      output csh4_clear_wr_t0_l                /* <ck1> */,
      output csh4_data_clr_done_l              /* <er2> */,
      output csh4_ebox_t0_in_h                 /* <fd1> */,
      output csh4_ebox_t3_l                    /* <au2> */,
      output csh4_ebox_wr_t4_in_h              /* <dh2> */,
      output csh4_one_word_wr_t0_l             /* <dj1> */,
      output csh4_writeback_t1_a_l             /* <fs1> */,
      output csh5_chan_rd_t5_l                 /* <ee2> */,
      output csh5_chan_t3_l                    /* <ad1> */,
      output csh5_chan_t4_l                    /* <ds2> */,
      output csh5_chan_wr_t5_in_h              /* <dr2> */,
      output csh5_page_refill_t12_l            /* <bt2> */,
      output csh5_page_refill_t4_l             /* <dj2> */,
      output csh5_page_refill_t8_l             /* <ar2> */,
      output csh5_page_refill_t9_l             /* <cj1> */,
      output csh5_t2_l                         /* <em1> */,
      output csh6_cache_wr_in_h                /* <am2> */,
      output csh6_cca_cyc_done_l               /* <dm2> */,
      output csh6_cca_inval_t4_l               /* <ap1> */,
      output csh6_chan_wr_cache_l              /* <ad2> */,
      output csh6_ebox_load_reg_h              /* <cn1> */,
      output csh6_mbox_pt_dir_wr_l             /* <cd2> */,
      output csh6_page_fail_hold_h             /* <cf2> */,
      output csh6_page_fail_hold_l             /* <df2> */,
      output csh6_page_refill_error_h          /* <bp1> */,
      output csh6_page_refill_error_l          /* <bm1> */,
      output csh6_wr_from_mem_nxt_h            /* <fp1> */,
      output csh7_cca_writeback_l              /* <el1> */,
      output csh7_e_writeback_l                /* <fk1> */,
      output csh7_fill_cache_rd_l              /* <ft2> */,
      input  csh_0_any_wr_l                    /* <ck2> */,
      input  csh_0_valid_match_h               /* <bj1> */,
      input  csh_0_valid_match_l               /* <cu2> */,
      input  csh_0_wd_val_h                    /* <de2> */,
      input  csh_1_any_wr_l                    /* <cm2> */,
      input  csh_1_valid_match_h               /* <bs2> */,
      input  csh_1_valid_match_l               /* <cv2> */,
      input  csh_1_wd_val_h                    /* <df1> */,
      input  csh_2_any_wr_l                    /* <cl2> */,
      input  csh_2_valid_match_h               /* <bv2> */,
      input  csh_2_valid_match_l               /* <ct2> */,
      input  csh_2_wd_val_h                    /* <dc1> */,
      input  csh_3_any_wr_l                    /* <cp1> */,
      input  csh_3_valid_match_h               /* <bs1> */,
      input  csh_3_valid_match_l               /* <cs2> */,
      input  csh_3_wd_val_h                    /* <dd2> */,
      output csh_chan_cyc_l                    /* <ak2> */,
      output csh_ebox_cyc_a_l                  /* <du2> */,
      input  csh_lru_1_h                       /* <cr1> */,
      input  csh_lru_2_h                       /* <cj2> */,
      output csh_refill_ram_wr_l               /* <fl2> */,
      output csh_use_hold_h                    /* <es2> */,
      output csh_use_wr_en_h                   /* <ar1> */,
      input  ctl3_diag_ld_ebus_reg_l           /* <dl2> */,
      input  diag_04_b_h                       /* <dp1> */,
      input  diag_05_b_h                       /* <dr1> */,
      input  diag_06_b_h                       /* <dm1> */,
      input  diag_read_func_17x_l              /* <ef1> */,
      output e_cache_wr_cyc_l                  /* <bh2> */,
      output ebus_d22_e_h                      /* <al1> */,
      output ebus_d23_e_h                      /* <am1> */,
      output ebus_d24_e_h                      /* <cd1> */,
      output ebus_d25_e_h                      /* <cm1> */,
      output ebus_d26_e_h                      /* <fd2> */,
      output ebus_d27_e_h                      /* <el2> */,
      output ebus_d28_e_h                      /* <er1> */,
      output ebus_d29_e_h                      /* <dk2> */,
      output load_ebus_reg_l                   /* <br1> */,
      output mb_test_par_a_in_l                /* <cf1> */,
      input  mbc1_write_ok_h                   /* <dd1> */,
      input  mbc2_csh_data_clr_t1_l            /* <af2> */,
      input  mbc2_csh_data_clr_t2_l            /* <bf1> */,
      input  mbc2_csh_data_clr_t3_l            /* <ek1> */,
      input  mbc2_data_clr_done_in_l           /* <eh2> */,
      input  mbc4_core_data_val_Ng1_l          /* <bl1> */,
      input  mbc4_core_data_valid_h            /* <ae1> */,
      input  mbc4_core_data_valid_l            /* <be1> */,
      input  mbx1_cache_bit_h                  /* <ah2> */,
      input  mbx1_cache_bit_l                  /* <ce2> */,
      input  mbx1_cca_all_pages_cyc_l          /* <bf2> */,
      input  mbx1_csh_cca_inval_csh_h          /* <al2> */,
      input  mbx1_csh_cca_val_core_h           /* <aj2> */,
      input  mbx1_csh_cca_val_core_l           /* <ac1> */,
      input  mbx1_refill_adr_en_nxt_h          /* <fc1> */,
      input  mbx2_mb_sel_hold_ff_h             /* <fu2> */,
      input  mbx2_mb_sel_hold_l                /* <cp2> */,
      input  mbx3_sbus_diag_3_l                /* <bd2> */,
      input  mbx4_cache_to_mb_done_l           /* <fk2> */,
      input  mbx5_mb_req_in_h                  /* <cs1> */,
      input  mcl2_vma_pause_h                  /* <ej1> */,
      input  mcl2_vma_read_l                   /* <fj2> */,
      input  mcl2_vma_write_l                  /* <dv2> */,
      input  mcl6_ebox_map_l                   /* <cl1> */,
      input  mem_busy_h                        /* <bl2> */,
      input  mr_reset_05_h                     /* <ae2> */,
      input  pag4_page_fail_l                  /* <as2> */,
      input  pag4_page_ok_l                    /* <ed1> */,
      input  pag4_page_refill_l                /* <dl1> */,
      input  phase_change_coming_l             /* <ed2> */,
      input  pma5_csh_writeback_cyc_l          /* <fp2> */,
      input  pma5_page_refill_cyc_l            /* <bm2> */,
      input  vma1_ac_ref_a_h                   /* <de1> */
);

`include "csh23nets.svh"

endmodule	// csh23
