// Triple 2 input XOR/XNOR
module mc10107(input bit a1, a2, b1, b2, c1, c2,
	       output bit qa, nqa,
	       output bit qb, nqb,
	       output bit qc, nqc);
  
  always_comb begin
    qa = a1 ^ a2;
    nqa = !qa;
    qb = b1 ^ b2;
    nqb = !qb;
    qc = c1 ^ c2;
    nqc = !qc;
  end
endmodule // mc10107
