// Framework for unit tests.

