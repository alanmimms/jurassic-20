module cra45(
      input  adEq0_l                           /* <da1> */,
      input  ad_00_h                           /* <ce2> */,
      input  ad_cry_Ng02_h                     /* <cf1> */,
      input  adx_00_a_h                        /* <dc1> */,
      input  ar_00_h                           /* <be2> */,
      input  ar_12_d_h                         /* <bu2> */,
      input  ar_18_d_h                         /* <cs2> */,
      input  arx_00_b_h                        /* <cv2> */,
      input  arx_01_b_h                        /* <dm1> */,
      input  arx_13_b_h                        /* <cs1> */,
      input  br_00_a_h                         /* <bv2> */,
      input  clk4_force_1777_h                 /* <bf2> */,
      input  clk4_pf_disp_07_h                 /* <ad1> */,
      input  clk4_pf_disp_08_h                 /* <ah2> */,
      input  clk4_pf_disp_09_h                 /* <ap1> */,
      input  clk4_pf_disp_10_h                 /* <bp2> */,
      input  clk_cra_h                         /* <cr2> */,
      input  con2_long_en_l                    /* <br2> */,
      input  con_cond_adr_10_h                 /* <de2> */,
      input  con_nicond_07_h                   /* <ac1> */,
      input  con_nicond_08_h                   /* <af2> */,
      input  con_nicond_09_h                   /* <am2> */,
      input  con_skip_en_40to47_l              /* <cr1> */,
      input  con_skip_en_50to57_l              /* <dd1> */,
      input  con_sr_00_h                       /* <ad2> */,
      input  con_sr_01_h                       /* <ak1> */,
      input  con_sr_02_h                       /* <an1> */,
      input  con_sr_03_h                       /* <bs1> */,
      input  cr02_dia_func_051_08_l            /* <ck1> */,
      input  cr02_dia_func_052_08_l            /* <ee1> */,
      input  cr02_dia_func_053_08_l            /* <at2> */,
      output cra1_adr_00_a_h                   /* <dl1> */,
      output cra1_adr_00_b_h                   /* <dp2> */,
      output cra1_adr_00_c_h                   /* <dk1> */,
      output cra1_adr_00_d_h                   /* <dj1> */,
      output cra1_adr_00_e_h                   /* <df2> */,
      output cra1_adr_01_a_l                   /* <fd1> */,
      output cra1_adr_01_b_h                   /* <fd2> */,
      output cra1_adr_01_c_l                   /* <fa1> */,
      output cra1_adr_01_d_h                   /* <fc1> */,
      output cra1_adr_01_e_l                   /* <et2> */,
      output cra1_adr_02_a_l                   /* <el1> */,
      output cra1_adr_02_b_h                   /* <ek1> */,
      output cra1_adr_02_c_l                   /* <el2> */,
      output cra1_adr_02_d_h                   /* <ek2> */,
      output cra1_adr_02_e_l                   /* <ef2> */,
      output cra1_adr_03_a_l                   /* <fp1> */,
      output cra1_adr_03_b_h                   /* <fs1> */,
      output cra1_adr_03_c_l                   /* <ft2> */,
      output cra1_adr_03_d_h                   /* <fr1> */,
      output cra1_adr_03_e_l                   /* <fn1> */,
      output cra1_adr_04_a_l                   /* <fl1> */,
      output cra1_adr_04_b_h                   /* <fl2> */,
      output cra1_adr_04_c_l                   /* <fh2> */,
      output cra1_adr_04_d_h                   /* <fk2> */,
      output cra1_adr_04_e_l                   /* <ff2> */,
      output cra1_adr_05_a_l                   /* <fr2> */,
      output cra1_adr_05_b_h                   /* <fu2> */,
      output cra1_adr_05_c_l                   /* <fp2> */,
      output cra1_adr_05_d_h                   /* <fs2> */,
      output cra1_adr_05_e_l                   /* <fm2> */,
      output cra1_adr_06_a_l                   /* <em1> */,
      output cra1_adr_06_b_h                   /* <ep1> */,
      output cra1_adr_06_c_l                   /* <en1> */,
      output cra1_adr_06_d_h                   /* <er1> */,
      output cra1_adr_06_e_l                   /* <ep2> */,
      output cra2_adr_07_a_h                   /* <cd1> */,
      output cra2_adr_07_b_h                   /* <ce1> */,
      output cra2_adr_07_c_h                   /* <cc1> */,
      output cra2_adr_07_d_h                   /* <cd2> */,
      output cra2_adr_07_e_h                   /* <ca1> */,
      output cra2_adr_08_a_h                   /* <au2> */,
      output cra2_adr_08_b_h                   /* <as2> */,
      output cra2_adr_08_c_h                   /* <ar2> */,
      output cra2_adr_08_d_h                   /* <ar1> */,
      output cra2_adr_08_e_h                   /* <as1> */,
      output cra2_adr_09_a_h                   /* <am1> */,
      output cra2_adr_09_b_h                   /* <al2> */,
      output cra2_adr_09_c_h                   /* <al1> */,
      output cra2_adr_09_d_h                   /* <ak2> */,
      output cra2_adr_09_e_h                   /* <aj2> */,
      output cra2_adr_10_a_h                   /* <ej1> */,
      output cra2_adr_10_b_h                   /* <ej2> */,
      output cra2_adr_10_c_h                   /* <eh2> */,
      output cra2_adr_10_d_h                   /* <ee2> */,
      output cra2_adr_10_e_h                   /* <ed2> */,
      input  cra2_spare_h                      /* <ct2> */,
      output cra3_disp_00_h                    /* <dm2> */,
      output cra3_disp_01_h                    /* <dt2> */,
      output cra3_disp_02_h                    /* <ef1> */,
      output cra3_disp_03_h                    /* <em2> */,
      output cra3_disp_04_h                    /* <es2> */,
      output cra3_disp_parity_h                /* <dl2> */,
      input  cram_cond_03s_h                   /* <cp2> */,
      input  cram_cond_04s_h                   /* <cp1> */,
      input  cram_cond_05s_h                   /* <cn1> */,
      input  cram_j00_h                        /* <dr2> */,
      input  cram_j01_h                        /* <fj1> */,
      input  cram_j02_h                        /* <fk1> */,
      input  cram_j03_h                        /* <fe2> */,
      input  cram_j04_h                        /* <fe1> */,
      input  cram_j05_h                        /* <be1> */,
      input  cram_j06_h                        /* <bd2> */,
      input  cram_j07_h                        /* <av2> */,
      input  cram_j08_h                        /* <ba1> */,
      input  cram_j09_h                        /* <ae2> */,
      input  cram_j10_h                        /* <af1> */,
      input  diag_04_a_l                       /* <dv2> */,
      input  diag_05_a_l                       /* <du2> */,
      input  diag_06_a_l                       /* <ds1> */,
      input  diag_read_func_14x_l              /* <bn1> */,
      input  dram_a_00_h                       /* <bm1> */,
      input  dram_a_01_h                       /* <bj2> */,
      input  dram_a_02_h                       /* <bk2> */,
      input  dram_b_00_h                       /* <bh2> */,
      input  dram_b_01_h                       /* <bl2> */,
      input  dram_b_02_h                       /* <cl1> */,
      input  dram_j_01_h                       /* <dp1> */,
      input  dram_j_02_h                       /* <dr1> */,
      input  dram_j_03_h                       /* <es1> */,
      input  dram_j_04_h                       /* <er2> */,
      input  dram_j_07_h                       /* <ae1> */,
      input  dram_j_08_h                       /* <bm2> */,
      input  dram_j_09_h                       /* <bj1> */,
      input  dram_j_10_h                       /* <bk1> */,
      input  ea_type_07_h                      /* <ff1> */,
      input  ea_type_08_h                      /* <ds2> */,
      input  ea_type_09_h                      /* <bs2> */,
      input  ea_type_10_h                      /* <cj2> */,
      output ebus_d00_e_h                      /* <dk2> */,
      output ebus_d01_e_h                      /* <dj2> */,
      output ebus_d02_e_h                      /* <df1> */,
      output ebus_d03_e_h                      /* <ed1> */,
      output ebus_d04_e_h                      /* <ec1> */,
      output ebus_d05_e_h                      /* <ea1> */,
      input  ir_acEq0_h                        /* <cm2> */,
      input  ir_norm_08_h                      /* <bd1> */,
      input  ir_norm_09_h                      /* <bt2> */,
      input  ir_norm_10_h                      /* <ck2> */,
      input  mcl6_pc_section_0_h               /* <dd2> */,
      input  mq_34_h                           /* <bl1> */,
      input  mq_35_h                           /* <cl2> */,
      input  mr_reset_04_h                     /* <dh2> */,
      input  scd1_scadEq0_l                    /* <de1> */,
      input  scd1_scad_sign_h                  /* <cf2> */,
      input  scd2_fe_sign_h                    /* <bf1> */,
      input  scd2_sc_sign_h                    /* <cm1> */,
      input  scd4_fpd_h                        /* <bc1> */,
      input  scd4_nicond_10_h                  /* <br1> */,
      input  shm1_ar_par_odd_b_l               /* <cu2> */,
      input  shm1_indexed_h                    /* <cj1> */,
      input  shm4_sh_00_a_h                    /* <aa1> */,
      input  shm4_sh_01_a_h                    /* <aj1> */,
      input  shm4_sh_02_a_h                    /* <ap2> */,
      input  shm4_sh_03_a_h                    /* <bp1> */,
      input  vma1_local_ac_address_l           /* <ch2> */
);

`include "cra45nets.svh"

endmodule	// cra45
