module tapped_delay_20_2(input bit in, output bit t1,t2,t3,t4,t5,t6,t7,t8,t9, out);
  always_comb t1 = in;
  always_comb t2 = in;
  always_comb t3 = in;
  always_comb t4 = in;
  always_comb t5 = in;
  always_comb t6 = in;
  always_comb t7 = in;
  always_comb t8 = in;
  always_comb t9 = in;
  always_comb out = in;
endmodule // tapped_delay_20_2
