module mb014(
  /* <fc1> */  input ar_12_a_h,
  /* <fd1> */  input ar_13_a_h,
  /* <eu2> */  input ar_14_a_h,
  /* <ev2> */  input ar_15_a_h,
  /* <cv2> */  input ar_16_a_h,
  /* <bu2> */  input ar_17_a_h,
  /* <dd2> */  input ar_30_a_h,
  /* <cs2> */  input ar_31_a_h,
  /* <bp1> */  input ar_32_a_h,
  /* <bj2> */  input ar_33_a_h,
  /* <bm2> */  input ar_34_a_h,
  /* <bf1> */  input ar_35_a_h,
  /* <er2> */  input cache_data_12_a_h,
  /* <ef1> */  input cache_data_13_a_h,
  /* <ff2> */  input cache_data_14_a_h,
  /* <er1> */  input cache_data_15_a_h,
  /* <cr1> */  input cache_data_16_a_h,
  /* <cm2> */  input cache_data_17_a_h,
  /* <dk2> */  input cache_data_30_a_h,
  /* <dk1> */  input cache_data_31_a_h,
  /* <am1> */  input cache_data_32_a_h,
  /* <ak1> */  input cache_data_33_a_h,
  /* <ar1> */  input cache_data_34_a_h,
  /* <ap1> */  input cache_data_35_a_h,
  /* <cj1> */  input cbus_d12_re_h,
  /* <ee1> */ output cbus_d12_te_h,
  /* <cj2> */  input cbus_d13_re_h,
  /* <ee2> */ output cbus_d13_te_h,
  /* <bs2> */  input cbus_d14_re_h,
  /* <el2> */ output cbus_d14_te_h,
  /* <bc1> */  input cbus_d15_re_h,
  /* <em1> */ output cbus_d15_te_h,
  /* <br1> */  input cbus_d16_re_h,
  /* <df1> */ output cbus_d16_te_h,
  /* <bd2> */  input cbus_d17_re_h,
  /* <dl2> */ output cbus_d17_te_h,
  /* <ch2> */  input cbus_d30_re_h,
  /* <dn1> */ output cbus_d30_te_h,
  /* <cf1> */  input cbus_d31_re_h,
  /* <dm2> */ output cbus_d31_te_h,
  /* <be2> */  input cbus_d32_re_h,
  /* <ah2> */ output cbus_d32_te_h,
  /* <bj1> */  input cbus_d33_re_h,
  /* <af2> */ output cbus_d33_te_h,
  /* <be1> */  input cbus_d34_re_h,
  /* <aj2> */ output cbus_d34_te_h,
  /* <bl1> */  input cbus_d35_re_h,
  /* <ak2> */ output cbus_d35_te_h,
  /* <fk1> */  input ccl_ccw_buf_wr_l,
  /* <ae2> */  input ccl_ch_buf_en_l,
  /* <es1> */  input ccl_mix_mb_sel_h,
  /* <fl1> */  input ccw_buf_12_in_h,
  /* <fm2> */  input ccw_buf_13_in_h,
  /* <fh2> */  input ccw_buf_14_in_h,
  /* <fj2> */  input ccw_buf_15_in_h,
  /* <cl2> */  input ccw_buf_16_in_h,
  /* <cl1> */  input ccw_buf_17_in_h,
  /* <ck2> */  input ccw_buf_30_in_h,
  /* <ck1> */  input ccw_buf_31_in_h,
  /* <at2> */  input ccw_buf_32_in_h,
  /* <as1> */  input ccw_buf_33_in_h,
  /* <ap2> */  input ccw_buf_34_in_h,
  /* <am2> */  input ccw_buf_35_in_h,
  /* <fk2> */  input ccw_buf_adr_0_h,
  /* <fj1> */  input ccw_buf_adr_1_h,
  /* <fl2> */  input ccw_buf_adr_2_h,
  /* <fm1> */  input ccw_buf_adr_3_h,
  /* <ek2> */ output ccw_mix_12_h,
  /* <eh2> */ output ccw_mix_13_h,
  /* <ff1> */ output ccw_mix_14_h,
  /* <es2> */ output ccw_mix_15_h,
  /* <cp2> */ output ccw_mix_16_h,
  /* <cn1> */ output ccw_mix_17_h,
  /* <dl1> */ output ccw_mix_30_h,
  /* <dh2> */ output ccw_mix_31_h,
  /* <al2> */ output ccw_mix_32_h,
  /* <al1> */ output ccw_mix_33_h,
  /* <as2> */ output ccw_mix_34_h,
  /* <ar2> */ output ccw_mix_35_h,
  /* <aj1> */  input ch_buf_wr_05_l,
  /* <ep1> */  input ch_buf_wr_2_l,
  /* <bd1> */  input ch_reverse_h,
  /* <fs2> */  input ch_t0_l,
  /* <af1> */  input ch_t2_l,
  /* <cr2> */  input clk_mb_12_h,
  /* <ek1> */  input con_ki10_paging_mode_l,
  /* <dt2> */  input crc_buf_mb_sel_h,
  /* <fu2> */  input crc_cbus_out_hold_h,
  /* <fp2> */  input crc_ch_buf_adr_0_h,
  /* <fr2> */  input crc_ch_buf_adr_1_h,
  /* <fp1> */  input crc_ch_buf_adr_2_h,
  /* <de1> */  input crc_ch_buf_adr_3_h,
  /* <dj1> */  input crc_ch_buf_adr_4_h,
  /* <de2> */  input crc_ch_buf_adr_5_h,
  /* <ae1> */  input crc_ch_buf_adr_6_h,
  /* <ad2> */  input mb0_hold_in_h,
  /* <ad1> */  input mb1_hold_in_h,
  /* <aa1> */  input mb2_hold_in_h,
  /* <ac1> */  input mb3_hold_in_h,
  /* <fc2> */  input mb_12_h,
  /* <fd2> */ output mb_12_h,
  /* <ds2> */ output mb_12to17_par_odd_h,
  /* <dr2> */ output mb_13_h,
  /* <dp2> */ output mb_14_h,
  /* <dm1> */ output mb_15_h,
  /* <dr1> */ output mb_16_h,
  /* <dp1> */ output mb_17_h,
  /* <av2> */ output mb_30_h,
  /* <au2> */ output mb_30to35_par_odd_h,
  /* <ba1> */ output mb_31_h,
  /* <cd2> */ output mb_32_h,
  /* <cd1> */ output mb_33_h,
  /* <ca1> */ output mb_34_h,
  /* <bv2> */ output mb_35_h,
  /* <ej1> */  input mb_in_sel_1_h,
  /* <el1> */  input mb_in_sel_2_h,
  /* <ep2> */  input mb_in_sel_4_h,
  /* <fr1> */  input mb_sel_1_en_h,
  /* <ft2> */  input mb_sel_2_en_h,
  /* <fv2> */  input mb_sel_hold_h,
  /* <em2> */  input mem_data_in_12_h,
  /* <ej2> */  input mem_data_in_13_h,
  /* <ea1> */  input mem_data_in_14_h,
  /* <dv2> */  input mem_data_in_15_h,
  /* <cp1> */  input mem_data_in_16_h,
  /* <cm1> */  input mem_data_in_17_h,
  /* <dj2> */  input mem_data_in_30_h,
  /* <df2> */  input mem_data_in_31_h,
  /* <bm1> */  input mem_data_in_32_h,
  /* <bk2> */  input mem_data_in_33_h,
  /* <bl2> */  input mem_data_in_34_h,
  /* <bk1> */  input mem_data_in_35_h,
  /* <ed2> */  input mem_to_c_en_l,
  /* <ed1> */  input mem_to_c_sel_1_h,
  /* <ds1> */  input mem_to_c_sel_2_h,
  /* <en1> */ output mem_to_cache_12_h,
  /* <ef2> */ output mem_to_cache_13_h,
  /* <ec1> */ output mem_to_cache_14_h,
  /* <du2> */ output mem_to_cache_15_h,
  /* <cf2> */ output mem_to_cache_16_h,
  /* <cc1> */ output mem_to_cache_17_h,
  /* <cs1> */ output mem_to_cache_30_h,
  /* <dd1> */ output mem_to_cache_31_h,
  /* <br2> */ output mem_to_cache_32_h,
  /* <bf2> */ output mem_to_cache_33_h,
  /* <bp2> */ output mem_to_cache_34_h,
  /* <bh2> */ output mem_to_cache_35_h,
  /* <fs1> */  input nxm_any_l,
  /* <fe1> */ output pt_in_12_h,
  /* <fe2> */ output pt_in_13_h,
  /* <fa1> */ output pt_in_14_h,
  /* <et2> */ output pt_in_15_h,
  /* <dc1> */ output pt_in_16_h,
  /* <da1> */ output pt_in_17_h,
  /* <cu2> */ output pt_in_30_h,
  /* <ct2> */ output pt_in_31_h,
  /* <ce1> */ output pt_in_32_h,
  /* <ce2> */ output pt_in_33_h,
  /* <bs1> */ output pt_in_34_h,
  /* <bt2> */ output pt_in_35_h
);

`include "mb014nets.svh"

endmodule	// mb014
