module ccw;
`include "ccw.svh"
endmodule	// ccw
