module mbx;
`include "mbx.svh"
endmodule	// mbx
