`ifndef __UTIL_SVH__
`define __UTIL_SVH__ 1

`define STRINGIFY(S)	`"S`"

`endif
