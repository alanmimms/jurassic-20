module chc09(
  /* <cl2> */  input cbus_ctom_e_h,
  /* <ds2> */  input cbus_done_e_h,
  /* <bh2> */ output cbus_error_e_h,
  /* <bf2> */ output cbus_last_word_e_h,
  /* <be2> */ output cbus_ready_e_h,
  /* <cs1> */  input cbus_request_e_h,
  /* <dv2> */  input cbus_reset_e_h,
  /* <ak1> */ output cbus_sel_0_e_h,
  /* <al1> */ output cbus_sel_1_e_h,
  /* <am1> */ output cbus_sel_2_e_h,
  /* <an1> */ output cbus_sel_3_e_h,
  /* <af1> */ output cbus_sel_4_e_h,
  /* <ae1> */ output cbus_sel_5_e_h,
  /* <ad1> */ output cbus_sel_6_e_h,
  /* <ac1> */ output cbus_sel_7_e_h,
  /* <dt2> */  input cbus_start_e_h,
  /* <du2> */  input cbus_store_e_h,
  /* <af2> */  input ccl_ch_buf_wr_en_l,
  /* <ch2> */  input ccl_mb_rip_l,
  /* <bs2> */  input ccw_diag_load_func_070_h,
  /* <el2> */ output ch_buf_wr_00_l,
  /* <em2> */ output ch_buf_wr_01_l,
  /* <ep2> */ output ch_buf_wr_02_l,
  /* <ek2> */ output ch_buf_wr_03_l,
  /* <ej2> */ output ch_buf_wr_04_l,
  /* <eh2> */ output ch_buf_wr_05_l,
  /* <br2> */ output ch_buf_wr_06_l,
  /* <at2> */ output ch_cbus_receive_ena_l,
  /* <bj2> */ output ch_cbus_req_h,
  /* <au2> */ output ch_cbus_req_l,
  /* <fm2> */ output ch_contr_1_l,
  /* <fp2> */ output ch_contr_2_l,
  /* <ft2> */ output ch_contr_4_l,
  /* <ce1> */ output ch_contr_req_h,
  /* <cf2> */ output ch_contr_req_l,
  /* <cd1> */ output ch_ctom_h,
  /* <bm2> */ output ch_ctom_l,
  /* <cc1> */ output ch_diag_04_h,
  /* <ak2> */ output ch_diag_04_l,
  /* <ca1> */ output ch_diag_05_h,
  /* <am2> */ output ch_diag_05_l,
  /* <aj1> */ output ch_diag_06_h,
  /* <fu2> */ output ch_diag_06_l,
  /* <ck2> */ output ch_diag_read_a_l,
  /* <as1> */ output ch_diag_read_b_l,
  /* <ar1> */ output ch_diag_read_c_l,
  /* <cs2> */ output ch_done_intr_h,
  /* <cu2> */ output ch_done_intr_l,
  /* <bu2> */ output ch_mb_req_inh_h,
  /* <bt2> */ output ch_mr_reset_b_h,
  /* <av2> */ output ch_req_d_l,
  /* <cp2> */ output ch_reset_intr_h,
  /* <fr2> */ output ch_reset_intr_l,
  /* <cf1> */ output ch_reverse_h,
  /* <ae2> */ output ch_sel_1b_en_l,
  /* <ad2> */ output ch_sel_2b_en_l,
  /* <ah2> */ output ch_sel_4b_en_l,
  /* <cm2> */ output ch_start_intr_h,
  /* <cv2> */ output ch_start_intr_l,
  /* <ef2> */ output ch_start_l,
  /* <cj2> */ output ch_store_h,
  /* <bk1> */ output ch_t0_h,
  /* <bp2> */ output ch_t0_l,
  /* <bl1> */ output ch_t1_h,
  /* <fv2> */ output ch_t1_l,
  /* <er2> */ output ch_t2_l,
  /* <bl2> */ output ch_t3_h,
  /* <aj2> */ output ch_t3_l,
  /* <as2> */ output chc1_cbus_out_ena_l,
  /* <bd2> */ output chc1_cbus_ready_e_l,
  /* <cr2> */  input clk1_chc_h,
  /* <ev2> */  input crc_cbus_contr_cyc_l,
  /* <dk2> */  input crc_err_in_h,
  /* <dr2> */  input crc_last_word_in_h,
  /* <ee2> */  input crc_ram_adr_1r_l,
  /* <ed2> */  input crc_ram_adr_2r_l,
  /* <ea1> */  input crc_ram_adr_4r_l,
  /* <dp2> */  input crc_ready_in_h,
  /* <dl2> */  input crc_reverse_in_h,
  /* <dd2> */  input crc_sel_1c_h,
  /* <es2> */  input crc_sel_1e_l,
  /* <df2> */  input crc_sel_2c_h,
  /* <et2> */  input crc_sel_2e_l,
  /* <de2> */  input crc_sel_4c_h,
  /* <eu2> */  input crc_sel_4e_l,
  /* <dm2> */  input crc_wr_ram_l,
  /* <al2> */  input diag_04_b_h,
  /* <ap2> */  input diag_05_b_h,
  /* <fs2> */  input diag_06_b_h,
  /* <ap1> */  input diag_read_func_17x_l,
  /* <bk2> */ output ebus_d00_e_h,
  /* <aa1> */ output ebus_d01_e_h,
  /* <bv2> */ output ebus_d02_e_h,
  /* <ce2> */ output ebus_d03_e_h,
  /* <df1> */  input ebus_d06_e_h,
  /* <dh2> */  input ebus_d07_e_h,
  /* <dj2> */  input ebus_d09_e_h,
  /* <dd1> */  input ebus_d10_e_h,
  /* <dc1> */  input ebus_d11_e_h,
  /* <da1> */  input ebus_d12_e_h,
  /* <ar2> */  input ebus_d13_e_h,
  /* <ct2> */  input mbc3_a_phase_coming_l,
  /* <cd2> */  input mr_reset_05_h
);

`include "chc09nets.svh"

endmodule	// chc09
