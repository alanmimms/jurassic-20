module mbc22(
      output a_change_coming_in_l              /* <ev2> */,
      output ackn_pulse_l                      /* <er1> */,
      input  apr2_wr_bad_adr_par_l             /* <es1> */,
      output cache_adr_27_h                    /* <aj2> */,
      output cache_adr_28_h                    /* <ak1> */,
      output cache_adr_29_h                    /* <ak2> */,
      output cache_adr_30_h                    /* <am2> */,
      output cache_adr_31_h                    /* <aa1> */,
      output cache_adr_32_h                    /* <ac1> */,
      output cache_adr_33_h                    /* <ad2> */,
      output cache_adr_34_h                    /* <cf1> */,
      output cache_adr_35_h                    /* <da1> */,
      output cache_adr_35_l                    /* <cm2> */,
      output cache_wr_00_a_l                   /* <cl2> */,
      output cache_wr_09_a_l                   /* <ck1> */,
      output cache_wr_18_a_l                   /* <ch2> */,
      output cache_wr_27_a_l                   /* <cj2> */,
      output cam_sel_1_h                       /* <cs2> */,
      output cam_sel_2_h                       /* <bj2> */,
      input  ccl_start_mem_l                   /* <df2> */,
      input  clk1_mbc_h                        /* <cr2> */,
      output core_busy_a_h                     /* <ee1> */,
      input  core_busy_h                       /* <ds1> */,
      output core_rd_in_prog_h                 /* <ef1> */,
      input  csh2_e_core_rd_rq_b_l             /* <dl2> */,
      input  csh2_one_word_rd_h                /* <et2> */,
      input  csh2_rd_pause_2nd_half_l          /* <el1> */,
      input  csh3_adr_pma_en_h                 /* <am1> */,
      input  csh3_any_val_hold_a_h             /* <df1> */,
      input  csh3_match_hold_1_in_h            /* <bf1> */,
      input  csh3_match_hold_2_in_h            /* <be2> */,
      output csh3_wr_en_l                      /* <cf2> */,
      input  csh4_clear_wr_t0_l                /* <dl1> */,
      input  csh4_data_clr_done_l              /* <es2> */,
      input  csh4_ebox_t3_l                    /* <dm2> */,
      input  csh4_ebox_wr_t4_in_h              /* <fn1> */,
      input  csh5_chan_rd_t5_l                 /* <cr1> */,
      input  csh5_chan_t3_l                    /* <dr1> */,
      input  csh5_chan_wr_t5_in_h              /* <fr2> */,
      input  csh5_page_refill_t9_l             /* <de1> */,
      input  csh6_cache_wr_in_h                /* <fl2> */,
      input  csh6_chan_wr_cache_l              /* <ep1> */,
      input  csh6_wr_from_mem_nxt_h            /* <fm2> */,
      output csh_0_wr_en_l                     /* <br1> */,
      output csh_1_wr_en_l                     /* <bd1> */,
      output csh_2_wr_en_l                     /* <dc1> */,
      output csh_adr_wr_pulse_l                /* <fl1> */,
      output csh_sel_lru_h                     /* <cp2> */,
      output csh_sel_lru_l                     /* <dm1> */,
      output csh_val_sel_all_h                 /* <cd2> */,
      output csh_val_wr_data_h                 /* <cn1> */,
      output csh_val_wr_pulse_l                /* <fp1> */,
      output csh_wr_sel_all_h                  /* <dj2> */,
      output csh_wr_wr_data_h                  /* <ek2> */,
      output csh_wr_wr_pulse_l                 /* <fp2> */,
      output data_valid_a_out_h                /* <br2> */,
      output data_valid_b_out_h                /* <dh2> */,
      input  diag_04_b_h                       /* <bc1> */,
      input  diag_05_b_h                       /* <ba1> */,
      input  diag_06_b_h                       /* <au2> */,
      input  diag_read_func_16x_l              /* <at2> */,
      input  e_cache_wr_cyc_l                  /* <eu2> */,
      output ebus_d27_e_h                      /* <cj1> */,
      output ebus_d28_e_h                      /* <cl1> */,
      output ebus_d29_e_h                      /* <ct2> */,
      output ebus_d30_e_h                      /* <dd1> */,
      output ebus_d31_e_h                      /* <dd2> */,
      output ebus_d32_e_h                      /* <dj1> */,
      output ebus_d33_e_h                      /* <dk1> */,
      output force_valid_match_0_h             /* <cu2> */,
      output force_valid_match_1_h             /* <bm1> */,
      output force_valid_match_2_h             /* <ca1> */,
      output force_valid_match_3_h             /* <cm1> */,
      input  load_ebus_reg_l                   /* <ae2> */,
      input  mb_sel_1_h                        /* <bs1> */,
      input  mb_sel_2_h                        /* <ce1> */,
      output mbc1_write_ok_h                   /* <ee2> */,
      output mbc2_csh_data_clr_t1_l            /* <cv2> */,
      output mbc2_csh_data_clr_t2_l            /* <bm2> */,
      output mbc2_csh_data_clr_t3_l            /* <cc1> */,
      output mbc2_data_clr_done_in_l           /* <bp2> */,
      output mbc3_a_change_coming_a_l          /* <ef2> */,
      output mbc3_a_phase_coming_l             /* <dk2> */,
      output mbc3_csh_wr_wr_data_l             /* <em2> */,
      output mbc3_inh_1st_mb_req_h             /* <bj1> */,
      output mbc4_core_adr_34_h                /* <ej2> */,
      output mbc4_core_adr_35_h                /* <bf2> */,
      output mbc4_core_data_val_Ng1_l          /* <bt2> */,
      output mbc4_core_data_val_Ng2_l          /* <ep2> */,
      output mbc4_core_data_valid_h            /* <ff2> */,
      output mbc4_core_data_valid_l            /* <fr1> */,
      output mbc4_mem_start_l                  /* <dv2> */,
      input  mbx1_cca_all_pages_cyc_l          /* <be1> */,
      input  mbx1_cca_inval_t4_a_h             /* <fm1> */,
      input  mbx1_force_match_en_l             /* <fa1> */,
      input  mbx1_refill_adr_en_h              /* <aj1> */,
      input  mbx2_chan_wr_cyc_l                /* <dp2> */,
      input  mbx3_refill_hold_h                /* <cd1> */,
      input  mbx4_cache_to_mb_t2_l             /* <em1> */,
      input  mbx4_cache_to_mb_t4_a_l           /* <dn1> */,
      input  mbx4_writeback_t2_h               /* <fs1> */,
      input  mbx5_mem_rd_rq_in_h               /* <fe1> */,
      input  mbx5_mem_to_c_en_l                /* <fc1> */,
      input  mbx5_mem_wr_rq_in_h               /* <fk1> */,
      input  mbx5_rq_0_in_h                    /* <fv2><fn2> */,
      input  mbx5_rq_1_in_h                    /* <fu2> */,
      input  mbx5_rq_2_in_h                    /* <ft2> */,
      input  mbx5_rq_3_in_h                    /* <fs2> */,
      output mbx_csh_adr_27_h                  /* <av2> */,
      output mbx_csh_adr_28_h                  /* <ap2> */,
      output mbx_csh_adr_29_h                  /* <ar2> */,
      output mbx_csh_adr_30_h                  /* <an1> */,
      output mbx_csh_adr_31_h                  /* <al1> */,
      output mbx_csh_adr_32_h                  /* <af2> */,
      output mbx_csh_adr_33_h                  /* <ad1> */,
      input  mem_ackn_a_h                      /* <ed2> */,
      input  mem_ackn_b_h                      /* <ed1> */,
      output mem_adr_par_h                     /* <bh2> */,
      input  mem_data_valid_a_l                /* <ea1> */,
      input  mem_data_valid_b_l                /* <ec1> */,
      output mem_rd_rq_b_h                     /* <cs1> */,
      output mem_rd_rq_h                       /* <ej1> */,
      output mem_rq_0_h                        /* <bk2> */,
      output mem_rq_1_h                        /* <bu2> */,
      output mem_rq_2_h                        /* <ck2> */,
      output mem_rq_3_h                        /* <du2> */,
      output mem_start_a_h                     /* <dr2> */,
      output mem_start_b_h                     /* <dp1> */,
      output mem_to_c_en_l                     /* <bs2> */,
      output mem_wr_rq_h                       /* <eh2> */,
      output mem_wr_rq_l                       /* <bl2> */,
      input  mr_reset_06_h                     /* <ce2> */,
      input  nxm_ackn_h                        /* <er2> */,
      input  nxm_data_val_l                    /* <fe2> */,
      output phase_change_coming_l             /* <en1> */,
      input  pma3_pa_27_h                      /* <bd2> */,
      input  pma3_pa_28_h                      /* <ar1> */,
      input  pma3_pa_29_h                      /* <as2> */,
      input  pma3_pa_30_h                      /* <af1> */,
      input  pma3_pa_31_h                      /* <al2> */,
      input  pma4_34_b_h                       /* <cp1> */,
      input  pma4_35_b_h                       /* <de2> */,
      input  pma4_adr_par_h                    /* <fk2> */,
      input  pma4_pa_32_h                      /* <ah2> */,
      input  pma4_pa_33_h                      /* <ae1> */,
      input  pma5_csh_writeback_cyc_l          /* <ds2> */,
      output rq_hold_ff_h                      /* <bp1> */,
      input  sbus_adr_34_h                     /* <fj2> */,
      input  sbus_adr_35_h                     /* <fj1> */,
      output sbus_adr_hold_h                   /* <dt2> */
);

`include "mbc22nets.svh"

endmodule	// mbc22
