module pic;
`include "pic.svh"
endmodule	// pic
